--------------------------------------------------------------------------------
-- Project      : Opallios
--------------------------------------------------------------------------------
-- File         : Opallios_FPGA_tb.vhd
-- Generated    : 07/06/2022
--------------------------------------------------------------------------------
-- Description  : Testbench for Opallios FPGA 
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library matrix;
use matrix.matrix_pkg.all;

entity Opallios_FPGA_tb is
end entity Opallios_FPGA_tb;

architecture rtl of Opallios_FPGA_tb is

    constant DEBUG : boolean := false;

    -- BeagleWire signals
    signal clk_100M    : std_logic;
    signal led         : std_logic_vector(3 downto 0);
    signal btn         : std_logic_vector(1 downto 0);
    signal sw          : std_logic_vector(1 downto 0);
    -- GPMC Interface
    signal gpmc_ad     : std_logic_vector(15 downto 0);
    signal gpmc_advn   : std_logic;
    signal gpmc_csn1   : std_logic;
    signal gpmc_wen    : std_logic;
    signal gpmc_oen    : std_logic;
    signal gpmc_clk    : std_logic;
    -- HUB75 interface
    signal R0          : std_logic;
    signal G0          : std_logic;
    signal B0          : std_logic;
    signal R1          : std_logic;
    signal G1          : std_logic;
    signal B1          : std_logic;
    signal Matrix_Addr : std_logic_vector(4 downto 0);
    signal Matrix_CLK  : std_logic;
    signal BLANK       : std_logic;
    signal LATCH       : std_logic;

    -- RGB Matrix array for TB
    signal MATRIX_TB   : t_RGB_matrix;

    -- Clock period definitions
    constant GPMC_CLK_period : time := 10 ns;

    component led_matrix_fpga_top is
        generic (
            DEBUG : boolean := false
        );
        port (
            -- BeagleWire signals
            clk_100M    : in  std_logic;
            led         : out std_logic_vector(3 downto 0);
            btn         : in  std_logic_vector(1 downto 0);
            sw          : in  std_logic_vector(1 downto 0);
            -- GPMC Interface
            gpmc_ad     : inout  std_logic_vector(15 downto 0);
            gpmc_advn   : in  std_logic;
            gpmc_csn1   : in  std_logic;
            gpmc_wen    : in  std_logic;
            gpmc_oen    : in  std_logic;
            gpmc_clk    : in  std_logic;
            -- HUB75 interface
            R0          : out std_logic;
            G0          : out std_logic;
            B0          : out std_logic;
            R1          : out std_logic;
            G1          : out std_logic;
            B1          : out std_logic;
            Matrix_Addr : out std_logic_vector(4 downto 0);
            Matrix_CLK  : out std_logic;
            BLANK       : out std_logic;
            LATCH       : out std_logic
        );
    end component;

    component matrix_64x64 is
    port (
        R0_IN       : in std_logic;
        G0_IN       : in std_logic;
        B0_IN       : in std_logic;
        R1_IN       : in std_logic;
        G1_IN       : in std_logic;
        B1_IN       : in std_logic;
        A_IN        : in std_logic_vector(4 downto 0);
        CLK_IN      : in std_logic;
        BLANK_IN    : in std_logic;
        LATCH_IN    : in std_logic;

        R0_OUT      : out std_logic;
        G0_OUT      : out std_logic;
        B0_OUT      : out std_logic;
        R1_OUT      : out std_logic;
        G1_OUT      : out std_logic;
        B1_OUT      : out std_logic;
        A_OUT       : out std_logic_vector(4 downto 0);
        CLK_OUT     : out std_logic;
        BLANK_OUT   : out std_logic;
        LATCH_OUT   : out std_logic;
        MATRIX_TB   : out t_RGB_matrix
    );
    end component;
        

begin

    --TB signals
    p_clk_100M : process
    begin
        clk_100M <= '1';
        wait for 5 ns;
        clk_100M <= '0';
        wait for 5 ns;
    end process;

    DUT: led_matrix_fpga_top
        generic map (
            DEBUG => DEBUG
        )
        port map (
            -- BeagleWire signals
            clk_100M    => clk_100M,
            led         => led,
            btn         => btn,
            sw          => sw,
            -- GPMC Interface
            gpmc_ad     => gpmc_ad,
            gpmc_advn   => gpmc_advn,
            gpmc_csn1   => gpmc_csn1,
            gpmc_wen    => gpmc_wen,
            gpmc_oen    => gpmc_oen,
            gpmc_clk    => gpmc_clk,
            -- HUB75 interface
            R0          => R0,
            G0          => G0,
            B0          => B0,
            R1          => R1,
            G1          => G1,
            B1          => B1,
            Matrix_Addr => Matrix_Addr,
            Matrix_CLK  => Matrix_CLK,
            BLANK       => BLANK,
            LATCH       => LATCH
        );

    u_matrix: matrix_64x64
        port map (
            R0_IN       => R0,
            G0_IN       => G0,
            B0_IN       => B0,
            R1_IN       => R1,
            G1_IN       => G1,
            B1_IN       => B1,
            A_IN        => Matrix_Addr,
            CLK_IN      => Matrix_CLK,
            BLANK_IN    => BLANK,
            LATCH_IN    => LATCH,

            R0_OUT      => open,
            G0_OUT      => open,
            B0_OUT      => open,
            R1_OUT      => open,
            G1_OUT      => open,
            B1_OUT      => open,
            A_OUT       => open,
            CLK_OUT     => open,
            BLANK_OUT   => open,
            LATCH_OUT   => open,
            MATRIX_TB   => MATRIX_TB
        );

    -- Clock process definitions
    p_GPMC_CLK :process
    begin
        GPMC_CLK <= '0';
        wait for GPMC_CLK_period/2;
        GPMC_CLK <= '1';
        wait for GPMC_CLK_period/2;
    end process;

    -- Stimulus process
    stim_proc: process
    procedure gpmc_send (RW   : std_logic;
                         ADDR : std_logic_vector(15 downto 0);
                         DATA : std_logic_vector(15 downto 0)) is
    begin
        
        GPMC_AD <= ADDR ;
        GPMC_CSN1 <= '0' ;
        GPMC_ADVN <= '0' ;
        GPMC_OEN <= '1' ;
        GPMC_WEN <= '1' ;
        wait for GPMC_CLK_period*2;
        GPMC_AD <= (others => 'Z') ;
        GPMC_CSN1 <= '0' ;
        GPMC_ADVN <= '1' ;
        GPMC_OEN <= '1' ;
        GPMC_WEN <= '1' ;
        wait for GPMC_CLK_period;
        if RW = '1' then 
            GPMC_AD <= DATA ;
            GPMC_CSN1 <= '0' ;
            GPMC_ADVN <= '1' ;
            GPMC_OEN <= '1' ;
            GPMC_WEN <= '0' ;     
        else 
            GPMC_AD <= (others => 'Z') ;
            GPMC_CSN1 <= '0' ;
            GPMC_ADVN <= '1' ;
            GPMC_OEN <= '0' ;
            GPMC_WEN <= '1' ;
        end if;
        wait for GPMC_CLK_period*4;
        GPMC_AD <= (others => 'Z') ;
        GPMC_CSN1 <= '1' ;
        GPMC_ADVN <= '1' ;
        GPMC_OEN <= '1' ;
        GPMC_WEN <= '1' ;
        wait for GPMC_CLK_period*10;
    end procedure gpmc_send;

    begin

        GPMC_AD <=  (others => 'Z');
        GPMC_CSN1 <= '1' ;
        GPMC_ADVN <= '1' ;
        GPMC_OEN <= '1' ;
        GPMC_WEN <= '1' ;

    -- wait for 100 ns;	
    -- wait for GPMC_CLK_period*2000;	
    wait for GPMC_CLK_period*10;
    -- gpmc_send format - RW: 0 read 1 write, ADDR, DATA
    -- read reg 0
    gpmc_send('0',x"0000",x"0000");
    -- write reg 0
    gpmc_send('1',x"0000",x"1234");
    -- read reg 0
    gpmc_send('0',x"0000",x"0000");
    -- read reg 1
    gpmc_send('0',x"0001",x"0000");
    -- read reg 0
    gpmc_send('0',x"0000",x"0000");

    -- Write some data to the video memory
    -- gpmc_send('1',x"2000",x"0FFF"); -- row 0 led 0
    -- gpmc_send('1',x"2001",x"003F"); -- row 0 led 0
    -- gpmc_send('1',x"2080",x"0FFF"); -- row 1 led 0
    -- gpmc_send('1',x"2081",x"003F"); -- row 1 led 0
    -- gpmc_send('1',x"20FE",x"0FFF"); -- row 1 led 63
    -- gpmc_send('1',x"20FF",x"003F"); -- row 1 led 63
    -- gpmc_send('1',x"2FFE",x"0FFF"); -- row 31 led 63
    -- gpmc_send('1',x"2FFF",x"003F"); -- row 31 led 63

    gpmc_send('1',x"2000",x"3F00");
    gpmc_send('1',x"2001",x"0000");
    gpmc_send('1',x"2002",x"3F01");
    gpmc_send('1',x"2003",x"0000");
    gpmc_send('1',x"2004",x"3E02");
    gpmc_send('1',x"2005",x"0000");
    gpmc_send('1',x"2006",x"3D03");
    gpmc_send('1',x"2007",x"0000");
    gpmc_send('1',x"2008",x"3C04");
    gpmc_send('1',x"2009",x"0000");
    gpmc_send('1',x"200A",x"3B05");
    gpmc_send('1',x"200B",x"0000");
    gpmc_send('1',x"200C",x"3A06");
    gpmc_send('1',x"200D",x"0000");
    gpmc_send('1',x"200E",x"3907");
    gpmc_send('1',x"200F",x"0000");
    gpmc_send('1',x"2010",x"3808");
    gpmc_send('1',x"2011",x"0000");
    gpmc_send('1',x"2012",x"3709");
    gpmc_send('1',x"2013",x"0000");
    gpmc_send('1',x"2014",x"360A");
    gpmc_send('1',x"2015",x"0000");
    gpmc_send('1',x"2016",x"350B");
    gpmc_send('1',x"2017",x"0000");
    gpmc_send('1',x"2018",x"340C");
    gpmc_send('1',x"2019",x"0000");
    gpmc_send('1',x"201A",x"330D");
    gpmc_send('1',x"201B",x"0000");
    gpmc_send('1',x"201C",x"320E");
    gpmc_send('1',x"201D",x"0000");
    gpmc_send('1',x"201E",x"310F");
    gpmc_send('1',x"201F",x"0000");
    gpmc_send('1',x"2020",x"3010");
    gpmc_send('1',x"2021",x"0000");
    gpmc_send('1',x"2022",x"2F11");
    gpmc_send('1',x"2023",x"0000");
    gpmc_send('1',x"2024",x"2E12");
    gpmc_send('1',x"2025",x"0000");
    gpmc_send('1',x"2026",x"2D13");
    gpmc_send('1',x"2027",x"0000");
    gpmc_send('1',x"2028",x"2C14");
    gpmc_send('1',x"2029",x"0000");
    gpmc_send('1',x"202A",x"2B15");
    gpmc_send('1',x"202B",x"0000");
    gpmc_send('1',x"202C",x"2A16");
    gpmc_send('1',x"202D",x"0000");
    gpmc_send('1',x"202E",x"2917");
    gpmc_send('1',x"202F",x"0000");
    gpmc_send('1',x"2030",x"2818");
    gpmc_send('1',x"2031",x"0000");
    gpmc_send('1',x"2032",x"2719");
    gpmc_send('1',x"2033",x"0000");
    gpmc_send('1',x"2034",x"261A");
    gpmc_send('1',x"2035",x"0000");
    gpmc_send('1',x"2036",x"251B");
    gpmc_send('1',x"2037",x"0000");
    gpmc_send('1',x"2038",x"241C");
    gpmc_send('1',x"2039",x"0000");
    gpmc_send('1',x"203A",x"231D");
    gpmc_send('1',x"203B",x"0000");
    gpmc_send('1',x"203C",x"221E");
    gpmc_send('1',x"203D",x"0000");
    gpmc_send('1',x"203E",x"211F");
    gpmc_send('1',x"203F",x"0000");
    gpmc_send('1',x"2040",x"2020");
    gpmc_send('1',x"2041",x"0000");
    gpmc_send('1',x"2042",x"1F21");
    gpmc_send('1',x"2043",x"0000");
    gpmc_send('1',x"2044",x"1E22");
    gpmc_send('1',x"2045",x"0000");
    gpmc_send('1',x"2046",x"1D23");
    gpmc_send('1',x"2047",x"0000");
    gpmc_send('1',x"2048",x"1C24");
    gpmc_send('1',x"2049",x"0000");
    gpmc_send('1',x"204A",x"1B25");
    gpmc_send('1',x"204B",x"0000");
    gpmc_send('1',x"204C",x"1A26");
    gpmc_send('1',x"204D",x"0000");
    gpmc_send('1',x"204E",x"1927");
    gpmc_send('1',x"204F",x"0000");
    gpmc_send('1',x"2050",x"1828");
    gpmc_send('1',x"2051",x"0000");
    gpmc_send('1',x"2052",x"1729");
    gpmc_send('1',x"2053",x"0000");
    gpmc_send('1',x"2054",x"162A");
    gpmc_send('1',x"2055",x"0000");
    gpmc_send('1',x"2056",x"152B");
    gpmc_send('1',x"2057",x"0000");
    gpmc_send('1',x"2058",x"142C");
    gpmc_send('1',x"2059",x"0000");
    gpmc_send('1',x"205A",x"132D");
    gpmc_send('1',x"205B",x"0000");
    gpmc_send('1',x"205C",x"122E");
    gpmc_send('1',x"205D",x"0000");
    gpmc_send('1',x"205E",x"112F");
    gpmc_send('1',x"205F",x"0000");
    gpmc_send('1',x"2060",x"1030");
    gpmc_send('1',x"2061",x"0000");
    gpmc_send('1',x"2062",x"0F31");
    gpmc_send('1',x"2063",x"0000");
    gpmc_send('1',x"2064",x"0E32");
    gpmc_send('1',x"2065",x"0000");
    gpmc_send('1',x"2066",x"0D33");
    gpmc_send('1',x"2067",x"0000");
    gpmc_send('1',x"2068",x"0C34");
    gpmc_send('1',x"2069",x"0000");
    gpmc_send('1',x"206A",x"0B35");
    gpmc_send('1',x"206B",x"0000");
    gpmc_send('1',x"206C",x"0A36");
    gpmc_send('1',x"206D",x"0000");
    gpmc_send('1',x"206E",x"0937");
    gpmc_send('1',x"206F",x"0000");
    gpmc_send('1',x"2070",x"0838");
    gpmc_send('1',x"2071",x"0000");
    gpmc_send('1',x"2072",x"0739");
    gpmc_send('1',x"2073",x"0000");
    gpmc_send('1',x"2074",x"063A");
    gpmc_send('1',x"2075",x"0000");
    gpmc_send('1',x"2076",x"053B");
    gpmc_send('1',x"2077",x"0000");
    gpmc_send('1',x"2078",x"043C");
    gpmc_send('1',x"2079",x"0000");
    gpmc_send('1',x"207A",x"033D");
    gpmc_send('1',x"207B",x"0000");
    gpmc_send('1',x"207C",x"023E");
    gpmc_send('1',x"207D",x"0000");
    gpmc_send('1',x"207E",x"013F");
    gpmc_send('1',x"207F",x"0000");
    gpmc_send('1',x"2080",x"003F");
    gpmc_send('1',x"2081",x"0000");
    gpmc_send('1',x"2082",x"003E");
    gpmc_send('1',x"2083",x"0001");
    gpmc_send('1',x"2084",x"003D");
    gpmc_send('1',x"2085",x"0002");
    gpmc_send('1',x"2086",x"003C");
    gpmc_send('1',x"2087",x"0003");
    gpmc_send('1',x"2088",x"003B");
    gpmc_send('1',x"2089",x"0004");
    gpmc_send('1',x"208A",x"003A");
    gpmc_send('1',x"208B",x"0005");
    gpmc_send('1',x"208C",x"0039");
    gpmc_send('1',x"208D",x"0006");
    gpmc_send('1',x"208E",x"0038");
    gpmc_send('1',x"208F",x"0007");
    gpmc_send('1',x"2090",x"0037");
    gpmc_send('1',x"2091",x"0008");
    gpmc_send('1',x"2092",x"0036");
    gpmc_send('1',x"2093",x"0009");
    gpmc_send('1',x"2094",x"0035");
    gpmc_send('1',x"2095",x"000A");
    gpmc_send('1',x"2096",x"0034");
    gpmc_send('1',x"2097",x"000B");
    gpmc_send('1',x"2098",x"0033");
    gpmc_send('1',x"2099",x"000C");
    gpmc_send('1',x"209A",x"0032");
    gpmc_send('1',x"209B",x"000D");
    gpmc_send('1',x"209C",x"0031");
    gpmc_send('1',x"209D",x"000E");
    gpmc_send('1',x"209E",x"0030");
    gpmc_send('1',x"209F",x"000F");
    gpmc_send('1',x"20A0",x"002F");
    gpmc_send('1',x"20A1",x"0010");
    gpmc_send('1',x"20A2",x"002E");
    gpmc_send('1',x"20A3",x"0011");
    gpmc_send('1',x"20A4",x"002D");
    gpmc_send('1',x"20A5",x"0012");
    gpmc_send('1',x"20A6",x"002C");
    gpmc_send('1',x"20A7",x"0013");
    gpmc_send('1',x"20A8",x"002B");
    gpmc_send('1',x"20A9",x"0014");
    gpmc_send('1',x"20AA",x"002A");
    gpmc_send('1',x"20AB",x"0015");
    gpmc_send('1',x"20AC",x"0029");
    gpmc_send('1',x"20AD",x"0016");
    gpmc_send('1',x"20AE",x"0028");
    gpmc_send('1',x"20AF",x"0017");
    gpmc_send('1',x"20B0",x"0027");
    gpmc_send('1',x"20B1",x"0018");
    gpmc_send('1',x"20B2",x"0026");
    gpmc_send('1',x"20B3",x"0019");
    gpmc_send('1',x"20B4",x"0025");
    gpmc_send('1',x"20B5",x"001A");
    gpmc_send('1',x"20B6",x"0024");
    gpmc_send('1',x"20B7",x"001B");
    gpmc_send('1',x"20B8",x"0023");
    gpmc_send('1',x"20B9",x"001C");
    gpmc_send('1',x"20BA",x"0022");
    gpmc_send('1',x"20BB",x"001D");
    gpmc_send('1',x"20BC",x"0021");
    gpmc_send('1',x"20BD",x"001E");
    gpmc_send('1',x"20BE",x"0020");
    gpmc_send('1',x"20BF",x"001F");
    gpmc_send('1',x"20C0",x"001F");
    gpmc_send('1',x"20C1",x"0020");
    gpmc_send('1',x"20C2",x"001E");
    gpmc_send('1',x"20C3",x"0021");
    gpmc_send('1',x"20C4",x"001D");
    gpmc_send('1',x"20C5",x"0022");
    gpmc_send('1',x"20C6",x"001C");
    gpmc_send('1',x"20C7",x"0023");
    gpmc_send('1',x"20C8",x"001B");
    gpmc_send('1',x"20C9",x"0024");
    gpmc_send('1',x"20CA",x"001A");
    gpmc_send('1',x"20CB",x"0025");
    gpmc_send('1',x"20CC",x"0019");
    gpmc_send('1',x"20CD",x"0026");
    gpmc_send('1',x"20CE",x"0018");
    gpmc_send('1',x"20CF",x"0027");
    gpmc_send('1',x"20D0",x"0017");
    gpmc_send('1',x"20D1",x"0028");
    gpmc_send('1',x"20D2",x"0016");
    gpmc_send('1',x"20D3",x"0029");
    gpmc_send('1',x"20D4",x"0015");
    gpmc_send('1',x"20D5",x"002A");
    gpmc_send('1',x"20D6",x"0014");
    gpmc_send('1',x"20D7",x"002B");
    gpmc_send('1',x"20D8",x"0013");
    gpmc_send('1',x"20D9",x"002C");
    gpmc_send('1',x"20DA",x"0012");
    gpmc_send('1',x"20DB",x"002D");
    gpmc_send('1',x"20DC",x"0011");
    gpmc_send('1',x"20DD",x"002E");
    gpmc_send('1',x"20DE",x"0010");
    gpmc_send('1',x"20DF",x"002F");
    gpmc_send('1',x"20E0",x"000F");
    gpmc_send('1',x"20E1",x"0030");
    gpmc_send('1',x"20E2",x"000E");
    gpmc_send('1',x"20E3",x"0031");
    gpmc_send('1',x"20E4",x"000D");
    gpmc_send('1',x"20E5",x"0032");
    gpmc_send('1',x"20E6",x"000C");
    gpmc_send('1',x"20E7",x"0033");
    gpmc_send('1',x"20E8",x"000B");
    gpmc_send('1',x"20E9",x"0034");
    gpmc_send('1',x"20EA",x"000A");
    gpmc_send('1',x"20EB",x"0035");
    gpmc_send('1',x"20EC",x"0009");
    gpmc_send('1',x"20ED",x"0036");
    gpmc_send('1',x"20EE",x"0008");
    gpmc_send('1',x"20EF",x"0037");
    gpmc_send('1',x"20F0",x"0007");
    gpmc_send('1',x"20F1",x"0038");
    gpmc_send('1',x"20F2",x"0006");
    gpmc_send('1',x"20F3",x"0039");
    gpmc_send('1',x"20F4",x"0005");
    gpmc_send('1',x"20F5",x"003A");
    gpmc_send('1',x"20F6",x"0004");
    gpmc_send('1',x"20F7",x"003B");
    gpmc_send('1',x"20F8",x"0003");
    gpmc_send('1',x"20F9",x"003C");
    gpmc_send('1',x"20FA",x"0002");
    gpmc_send('1',x"20FB",x"003D");
    gpmc_send('1',x"20FC",x"0001");
    gpmc_send('1',x"20FD",x"003E");
    gpmc_send('1',x"20FE",x"0000");
    gpmc_send('1',x"20FF",x"003F");
    gpmc_send('1',x"2100",x"0100");
    gpmc_send('1',x"2101",x"003E");
    gpmc_send('1',x"2102",x"0200");
    gpmc_send('1',x"2103",x"003D");
    gpmc_send('1',x"2104",x"0300");
    gpmc_send('1',x"2105",x"003C");
    gpmc_send('1',x"2106",x"0400");
    gpmc_send('1',x"2107",x"003B");
    gpmc_send('1',x"2108",x"0500");
    gpmc_send('1',x"2109",x"003A");
    gpmc_send('1',x"210A",x"0600");
    gpmc_send('1',x"210B",x"0039");
    gpmc_send('1',x"210C",x"0700");
    gpmc_send('1',x"210D",x"0038");
    gpmc_send('1',x"210E",x"0800");
    gpmc_send('1',x"210F",x"0037");
    gpmc_send('1',x"2110",x"0900");
    gpmc_send('1',x"2111",x"0036");
    gpmc_send('1',x"2112",x"0A00");
    gpmc_send('1',x"2113",x"0035");
    gpmc_send('1',x"2114",x"0B00");
    gpmc_send('1',x"2115",x"0034");
    gpmc_send('1',x"2116",x"0C00");
    gpmc_send('1',x"2117",x"0033");
    gpmc_send('1',x"2118",x"0D00");
    gpmc_send('1',x"2119",x"0032");
    gpmc_send('1',x"211A",x"0E00");
    gpmc_send('1',x"211B",x"0031");
    gpmc_send('1',x"211C",x"0F00");
    gpmc_send('1',x"211D",x"0030");
    gpmc_send('1',x"211E",x"1000");
    gpmc_send('1',x"211F",x"002F");
    gpmc_send('1',x"2120",x"1100");
    gpmc_send('1',x"2121",x"002E");
    gpmc_send('1',x"2122",x"1200");
    gpmc_send('1',x"2123",x"002D");
    gpmc_send('1',x"2124",x"1300");
    gpmc_send('1',x"2125",x"002C");
    gpmc_send('1',x"2126",x"1400");
    gpmc_send('1',x"2127",x"002B");
    gpmc_send('1',x"2128",x"1500");
    gpmc_send('1',x"2129",x"002A");
    gpmc_send('1',x"212A",x"1600");
    gpmc_send('1',x"212B",x"0029");
    gpmc_send('1',x"212C",x"1700");
    gpmc_send('1',x"212D",x"0028");
    gpmc_send('1',x"212E",x"1800");
    gpmc_send('1',x"212F",x"0027");
    gpmc_send('1',x"2130",x"1900");
    gpmc_send('1',x"2131",x"0026");
    gpmc_send('1',x"2132",x"1A00");
    gpmc_send('1',x"2133",x"0025");
    gpmc_send('1',x"2134",x"1B00");
    gpmc_send('1',x"2135",x"0024");
    gpmc_send('1',x"2136",x"1C00");
    gpmc_send('1',x"2137",x"0023");
    gpmc_send('1',x"2138",x"1D00");
    gpmc_send('1',x"2139",x"0022");
    gpmc_send('1',x"213A",x"1E00");
    gpmc_send('1',x"213B",x"0021");
    gpmc_send('1',x"213C",x"1F00");
    gpmc_send('1',x"213D",x"0020");
    gpmc_send('1',x"213E",x"2000");
    gpmc_send('1',x"213F",x"001F");
    gpmc_send('1',x"2140",x"2100");
    gpmc_send('1',x"2141",x"001E");
    gpmc_send('1',x"2142",x"2200");
    gpmc_send('1',x"2143",x"001D");
    gpmc_send('1',x"2144",x"2300");
    gpmc_send('1',x"2145",x"001C");
    gpmc_send('1',x"2146",x"2400");
    gpmc_send('1',x"2147",x"001B");
    gpmc_send('1',x"2148",x"2500");
    gpmc_send('1',x"2149",x"001A");
    gpmc_send('1',x"214A",x"2600");
    gpmc_send('1',x"214B",x"0019");
    gpmc_send('1',x"214C",x"2700");
    gpmc_send('1',x"214D",x"0018");
    gpmc_send('1',x"214E",x"2800");
    gpmc_send('1',x"214F",x"0017");
    gpmc_send('1',x"2150",x"2900");
    gpmc_send('1',x"2151",x"0016");
    gpmc_send('1',x"2152",x"2A00");
    gpmc_send('1',x"2153",x"0015");
    gpmc_send('1',x"2154",x"2B00");
    gpmc_send('1',x"2155",x"0014");
    gpmc_send('1',x"2156",x"2C00");
    gpmc_send('1',x"2157",x"0013");
    gpmc_send('1',x"2158",x"2D00");
    gpmc_send('1',x"2159",x"0012");
    gpmc_send('1',x"215A",x"2E00");
    gpmc_send('1',x"215B",x"0011");
    gpmc_send('1',x"215C",x"2F00");
    gpmc_send('1',x"215D",x"0010");
    gpmc_send('1',x"215E",x"3000");
    gpmc_send('1',x"215F",x"000F");
    gpmc_send('1',x"2160",x"3100");
    gpmc_send('1',x"2161",x"000E");
    gpmc_send('1',x"2162",x"3200");
    gpmc_send('1',x"2163",x"000D");
    gpmc_send('1',x"2164",x"3300");
    gpmc_send('1',x"2165",x"000C");
    gpmc_send('1',x"2166",x"3400");
    gpmc_send('1',x"2167",x"000B");
    gpmc_send('1',x"2168",x"3500");
    gpmc_send('1',x"2169",x"000A");
    gpmc_send('1',x"216A",x"3600");
    gpmc_send('1',x"216B",x"0009");
    gpmc_send('1',x"216C",x"3700");
    gpmc_send('1',x"216D",x"0008");
    gpmc_send('1',x"216E",x"3800");
    gpmc_send('1',x"216F",x"0007");
    gpmc_send('1',x"2170",x"3900");
    gpmc_send('1',x"2171",x"0006");
    gpmc_send('1',x"2172",x"3A00");
    gpmc_send('1',x"2173",x"0005");
    gpmc_send('1',x"2174",x"3B00");
    gpmc_send('1',x"2175",x"0004");
    gpmc_send('1',x"2176",x"3C00");
    gpmc_send('1',x"2177",x"0003");
    gpmc_send('1',x"2178",x"3D00");
    gpmc_send('1',x"2179",x"0002");
    gpmc_send('1',x"217A",x"3E00");
    gpmc_send('1',x"217B",x"0001");
    gpmc_send('1',x"217C",x"3F00");
    gpmc_send('1',x"217D",x"0000");
    gpmc_send('1',x"217E",x"3F01");
    gpmc_send('1',x"217F",x"0000");
    gpmc_send('1',x"2180",x"3E02");
    gpmc_send('1',x"2181",x"0000");
    gpmc_send('1',x"2182",x"3D03");
    gpmc_send('1',x"2183",x"0000");
    gpmc_send('1',x"2184",x"3C04");
    gpmc_send('1',x"2185",x"0000");
    gpmc_send('1',x"2186",x"3B05");
    gpmc_send('1',x"2187",x"0000");
    gpmc_send('1',x"2188",x"3A06");
    gpmc_send('1',x"2189",x"0000");
    gpmc_send('1',x"218A",x"3907");
    gpmc_send('1',x"218B",x"0000");
    gpmc_send('1',x"218C",x"3808");
    gpmc_send('1',x"218D",x"0000");
    gpmc_send('1',x"218E",x"3709");
    gpmc_send('1',x"218F",x"0000");
    gpmc_send('1',x"2190",x"360A");
    gpmc_send('1',x"2191",x"0000");
    gpmc_send('1',x"2192",x"350B");
    gpmc_send('1',x"2193",x"0000");
    gpmc_send('1',x"2194",x"340C");
    gpmc_send('1',x"2195",x"0000");
    gpmc_send('1',x"2196",x"330D");
    gpmc_send('1',x"2197",x"0000");
    gpmc_send('1',x"2198",x"320E");
    gpmc_send('1',x"2199",x"0000");
    gpmc_send('1',x"219A",x"310F");
    gpmc_send('1',x"219B",x"0000");
    gpmc_send('1',x"219C",x"3010");
    gpmc_send('1',x"219D",x"0000");
    gpmc_send('1',x"219E",x"2F11");
    gpmc_send('1',x"219F",x"0000");
    gpmc_send('1',x"21A0",x"2E12");
    gpmc_send('1',x"21A1",x"0000");
    gpmc_send('1',x"21A2",x"2D13");
    gpmc_send('1',x"21A3",x"0000");
    gpmc_send('1',x"21A4",x"2C14");
    gpmc_send('1',x"21A5",x"0000");
    gpmc_send('1',x"21A6",x"2B15");
    gpmc_send('1',x"21A7",x"0000");
    gpmc_send('1',x"21A8",x"2A16");
    gpmc_send('1',x"21A9",x"0000");
    gpmc_send('1',x"21AA",x"2917");
    gpmc_send('1',x"21AB",x"0000");
    gpmc_send('1',x"21AC",x"2818");
    gpmc_send('1',x"21AD",x"0000");
    gpmc_send('1',x"21AE",x"2719");
    gpmc_send('1',x"21AF",x"0000");
    gpmc_send('1',x"21B0",x"261A");
    gpmc_send('1',x"21B1",x"0000");
    gpmc_send('1',x"21B2",x"251B");
    gpmc_send('1',x"21B3",x"0000");
    gpmc_send('1',x"21B4",x"241C");
    gpmc_send('1',x"21B5",x"0000");
    gpmc_send('1',x"21B6",x"231D");
    gpmc_send('1',x"21B7",x"0000");
    gpmc_send('1',x"21B8",x"221E");
    gpmc_send('1',x"21B9",x"0000");
    gpmc_send('1',x"21BA",x"211F");
    gpmc_send('1',x"21BB",x"0000");
    gpmc_send('1',x"21BC",x"2020");
    gpmc_send('1',x"21BD",x"0000");
    gpmc_send('1',x"21BE",x"1F21");
    gpmc_send('1',x"21BF",x"0000");
    gpmc_send('1',x"21C0",x"1E22");
    gpmc_send('1',x"21C1",x"0000");
    gpmc_send('1',x"21C2",x"1D23");
    gpmc_send('1',x"21C3",x"0000");
    gpmc_send('1',x"21C4",x"1C24");
    gpmc_send('1',x"21C5",x"0000");
    gpmc_send('1',x"21C6",x"1B25");
    gpmc_send('1',x"21C7",x"0000");
    gpmc_send('1',x"21C8",x"1A26");
    gpmc_send('1',x"21C9",x"0000");
    gpmc_send('1',x"21CA",x"1927");
    gpmc_send('1',x"21CB",x"0000");
    gpmc_send('1',x"21CC",x"1828");
    gpmc_send('1',x"21CD",x"0000");
    gpmc_send('1',x"21CE",x"1729");
    gpmc_send('1',x"21CF",x"0000");
    gpmc_send('1',x"21D0",x"162A");
    gpmc_send('1',x"21D1",x"0000");
    gpmc_send('1',x"21D2",x"152B");
    gpmc_send('1',x"21D3",x"0000");
    gpmc_send('1',x"21D4",x"142C");
    gpmc_send('1',x"21D5",x"0000");
    gpmc_send('1',x"21D6",x"132D");
    gpmc_send('1',x"21D7",x"0000");
    gpmc_send('1',x"21D8",x"122E");
    gpmc_send('1',x"21D9",x"0000");
    gpmc_send('1',x"21DA",x"112F");
    gpmc_send('1',x"21DB",x"0000");
    gpmc_send('1',x"21DC",x"1030");
    gpmc_send('1',x"21DD",x"0000");
    gpmc_send('1',x"21DE",x"0F31");
    gpmc_send('1',x"21DF",x"0000");
    gpmc_send('1',x"21E0",x"0E32");
    gpmc_send('1',x"21E1",x"0000");
    gpmc_send('1',x"21E2",x"0D33");
    gpmc_send('1',x"21E3",x"0000");
    gpmc_send('1',x"21E4",x"0C34");
    gpmc_send('1',x"21E5",x"0000");
    gpmc_send('1',x"21E6",x"0B35");
    gpmc_send('1',x"21E7",x"0000");
    gpmc_send('1',x"21E8",x"0A36");
    gpmc_send('1',x"21E9",x"0000");
    gpmc_send('1',x"21EA",x"0937");
    gpmc_send('1',x"21EB",x"0000");
    gpmc_send('1',x"21EC",x"0838");
    gpmc_send('1',x"21ED",x"0000");
    gpmc_send('1',x"21EE",x"0739");
    gpmc_send('1',x"21EF",x"0000");
    gpmc_send('1',x"21F0",x"063A");
    gpmc_send('1',x"21F1",x"0000");
    gpmc_send('1',x"21F2",x"053B");
    gpmc_send('1',x"21F3",x"0000");
    gpmc_send('1',x"21F4",x"043C");
    gpmc_send('1',x"21F5",x"0000");
    gpmc_send('1',x"21F6",x"033D");
    gpmc_send('1',x"21F7",x"0000");
    gpmc_send('1',x"21F8",x"023E");
    gpmc_send('1',x"21F9",x"0000");
    gpmc_send('1',x"21FA",x"013F");
    gpmc_send('1',x"21FB",x"0000");
    gpmc_send('1',x"21FC",x"003F");
    gpmc_send('1',x"21FD",x"0000");
    gpmc_send('1',x"21FE",x"003E");
    gpmc_send('1',x"21FF",x"0001");
    gpmc_send('1',x"2200",x"003D");
    gpmc_send('1',x"2201",x"0002");
    gpmc_send('1',x"2202",x"003C");
    gpmc_send('1',x"2203",x"0003");
    gpmc_send('1',x"2204",x"003B");
    gpmc_send('1',x"2205",x"0004");
    gpmc_send('1',x"2206",x"003A");
    gpmc_send('1',x"2207",x"0005");
    gpmc_send('1',x"2208",x"0039");
    gpmc_send('1',x"2209",x"0006");
    gpmc_send('1',x"220A",x"0038");
    gpmc_send('1',x"220B",x"0007");
    gpmc_send('1',x"220C",x"0037");
    gpmc_send('1',x"220D",x"0008");
    gpmc_send('1',x"220E",x"0036");
    gpmc_send('1',x"220F",x"0009");
    gpmc_send('1',x"2210",x"0035");
    gpmc_send('1',x"2211",x"000A");
    gpmc_send('1',x"2212",x"0034");
    gpmc_send('1',x"2213",x"000B");
    gpmc_send('1',x"2214",x"0033");
    gpmc_send('1',x"2215",x"000C");
    gpmc_send('1',x"2216",x"0032");
    gpmc_send('1',x"2217",x"000D");
    gpmc_send('1',x"2218",x"0031");
    gpmc_send('1',x"2219",x"000E");
    gpmc_send('1',x"221A",x"0030");
    gpmc_send('1',x"221B",x"000F");
    gpmc_send('1',x"221C",x"002F");
    gpmc_send('1',x"221D",x"0010");
    gpmc_send('1',x"221E",x"002E");
    gpmc_send('1',x"221F",x"0011");
    gpmc_send('1',x"2220",x"002D");
    gpmc_send('1',x"2221",x"0012");
    gpmc_send('1',x"2222",x"002C");
    gpmc_send('1',x"2223",x"0013");
    gpmc_send('1',x"2224",x"002B");
    gpmc_send('1',x"2225",x"0014");
    gpmc_send('1',x"2226",x"002A");
    gpmc_send('1',x"2227",x"0015");
    gpmc_send('1',x"2228",x"0029");
    gpmc_send('1',x"2229",x"0016");
    gpmc_send('1',x"222A",x"0028");
    gpmc_send('1',x"222B",x"0017");
    gpmc_send('1',x"222C",x"0027");
    gpmc_send('1',x"222D",x"0018");
    gpmc_send('1',x"222E",x"0026");
    gpmc_send('1',x"222F",x"0019");
    gpmc_send('1',x"2230",x"0025");
    gpmc_send('1',x"2231",x"001A");
    gpmc_send('1',x"2232",x"0024");
    gpmc_send('1',x"2233",x"001B");
    gpmc_send('1',x"2234",x"0023");
    gpmc_send('1',x"2235",x"001C");
    gpmc_send('1',x"2236",x"0022");
    gpmc_send('1',x"2237",x"001D");
    gpmc_send('1',x"2238",x"0021");
    gpmc_send('1',x"2239",x"001E");
    gpmc_send('1',x"223A",x"0020");
    gpmc_send('1',x"223B",x"001F");
    gpmc_send('1',x"223C",x"001F");
    gpmc_send('1',x"223D",x"0020");
    gpmc_send('1',x"223E",x"001E");
    gpmc_send('1',x"223F",x"0021");
    gpmc_send('1',x"2240",x"001D");
    gpmc_send('1',x"2241",x"0022");
    gpmc_send('1',x"2242",x"001C");
    gpmc_send('1',x"2243",x"0023");
    gpmc_send('1',x"2244",x"001B");
    gpmc_send('1',x"2245",x"0024");
    gpmc_send('1',x"2246",x"001A");
    gpmc_send('1',x"2247",x"0025");
    gpmc_send('1',x"2248",x"0019");
    gpmc_send('1',x"2249",x"0026");
    gpmc_send('1',x"224A",x"0018");
    gpmc_send('1',x"224B",x"0027");
    gpmc_send('1',x"224C",x"0017");
    gpmc_send('1',x"224D",x"0028");
    gpmc_send('1',x"224E",x"0016");
    gpmc_send('1',x"224F",x"0029");
    gpmc_send('1',x"2250",x"0015");
    gpmc_send('1',x"2251",x"002A");
    gpmc_send('1',x"2252",x"0014");
    gpmc_send('1',x"2253",x"002B");
    gpmc_send('1',x"2254",x"0013");
    gpmc_send('1',x"2255",x"002C");
    gpmc_send('1',x"2256",x"0012");
    gpmc_send('1',x"2257",x"002D");
    gpmc_send('1',x"2258",x"0011");
    gpmc_send('1',x"2259",x"002E");
    gpmc_send('1',x"225A",x"0010");
    gpmc_send('1',x"225B",x"002F");
    gpmc_send('1',x"225C",x"000F");
    gpmc_send('1',x"225D",x"0030");
    gpmc_send('1',x"225E",x"000E");
    gpmc_send('1',x"225F",x"0031");
    gpmc_send('1',x"2260",x"000D");
    gpmc_send('1',x"2261",x"0032");
    gpmc_send('1',x"2262",x"000C");
    gpmc_send('1',x"2263",x"0033");
    gpmc_send('1',x"2264",x"000B");
    gpmc_send('1',x"2265",x"0034");
    gpmc_send('1',x"2266",x"000A");
    gpmc_send('1',x"2267",x"0035");
    gpmc_send('1',x"2268",x"0009");
    gpmc_send('1',x"2269",x"0036");
    gpmc_send('1',x"226A",x"0008");
    gpmc_send('1',x"226B",x"0037");
    gpmc_send('1',x"226C",x"0007");
    gpmc_send('1',x"226D",x"0038");
    gpmc_send('1',x"226E",x"0006");
    gpmc_send('1',x"226F",x"0039");
    gpmc_send('1',x"2270",x"0005");
    gpmc_send('1',x"2271",x"003A");
    gpmc_send('1',x"2272",x"0004");
    gpmc_send('1',x"2273",x"003B");
    gpmc_send('1',x"2274",x"0003");
    gpmc_send('1',x"2275",x"003C");
    gpmc_send('1',x"2276",x"0002");
    gpmc_send('1',x"2277",x"003D");
    gpmc_send('1',x"2278",x"0001");
    gpmc_send('1',x"2279",x"003E");
    gpmc_send('1',x"227A",x"0000");
    gpmc_send('1',x"227B",x"003F");
    gpmc_send('1',x"227C",x"0100");
    gpmc_send('1',x"227D",x"003E");
    gpmc_send('1',x"227E",x"0200");
    gpmc_send('1',x"227F",x"003D");
    gpmc_send('1',x"2280",x"0300");
    gpmc_send('1',x"2281",x"003C");
    gpmc_send('1',x"2282",x"0400");
    gpmc_send('1',x"2283",x"003B");
    gpmc_send('1',x"2284",x"0500");
    gpmc_send('1',x"2285",x"003A");
    gpmc_send('1',x"2286",x"0600");
    gpmc_send('1',x"2287",x"0039");
    gpmc_send('1',x"2288",x"0700");
    gpmc_send('1',x"2289",x"0038");
    gpmc_send('1',x"228A",x"0800");
    gpmc_send('1',x"228B",x"0037");
    gpmc_send('1',x"228C",x"0900");
    gpmc_send('1',x"228D",x"0036");
    gpmc_send('1',x"228E",x"0A00");
    gpmc_send('1',x"228F",x"0035");
    gpmc_send('1',x"2290",x"0B00");
    gpmc_send('1',x"2291",x"0034");
    gpmc_send('1',x"2292",x"0C00");
    gpmc_send('1',x"2293",x"0033");
    gpmc_send('1',x"2294",x"0D00");
    gpmc_send('1',x"2295",x"0032");
    gpmc_send('1',x"2296",x"0E00");
    gpmc_send('1',x"2297",x"0031");
    gpmc_send('1',x"2298",x"0F00");
    gpmc_send('1',x"2299",x"0030");
    gpmc_send('1',x"229A",x"1000");
    gpmc_send('1',x"229B",x"002F");
    gpmc_send('1',x"229C",x"1100");
    gpmc_send('1',x"229D",x"002E");
    gpmc_send('1',x"229E",x"1200");
    gpmc_send('1',x"229F",x"002D");
    gpmc_send('1',x"22A0",x"1300");
    gpmc_send('1',x"22A1",x"002C");
    gpmc_send('1',x"22A2",x"1400");
    gpmc_send('1',x"22A3",x"002B");
    gpmc_send('1',x"22A4",x"1500");
    gpmc_send('1',x"22A5",x"002A");
    gpmc_send('1',x"22A6",x"1600");
    gpmc_send('1',x"22A7",x"0029");
    gpmc_send('1',x"22A8",x"1700");
    gpmc_send('1',x"22A9",x"0028");
    gpmc_send('1',x"22AA",x"1800");
    gpmc_send('1',x"22AB",x"0027");
    gpmc_send('1',x"22AC",x"1900");
    gpmc_send('1',x"22AD",x"0026");
    gpmc_send('1',x"22AE",x"1A00");
    gpmc_send('1',x"22AF",x"0025");
    gpmc_send('1',x"22B0",x"1B00");
    gpmc_send('1',x"22B1",x"0024");
    gpmc_send('1',x"22B2",x"1C00");
    gpmc_send('1',x"22B3",x"0023");
    gpmc_send('1',x"22B4",x"1D00");
    gpmc_send('1',x"22B5",x"0022");
    gpmc_send('1',x"22B6",x"1E00");
    gpmc_send('1',x"22B7",x"0021");
    gpmc_send('1',x"22B8",x"1F00");
    gpmc_send('1',x"22B9",x"0020");
    gpmc_send('1',x"22BA",x"2000");
    gpmc_send('1',x"22BB",x"001F");
    gpmc_send('1',x"22BC",x"2100");
    gpmc_send('1',x"22BD",x"001E");
    gpmc_send('1',x"22BE",x"2200");
    gpmc_send('1',x"22BF",x"001D");
    gpmc_send('1',x"22C0",x"2300");
    gpmc_send('1',x"22C1",x"001C");
    gpmc_send('1',x"22C2",x"2400");
    gpmc_send('1',x"22C3",x"001B");
    gpmc_send('1',x"22C4",x"2500");
    gpmc_send('1',x"22C5",x"001A");
    gpmc_send('1',x"22C6",x"2600");
    gpmc_send('1',x"22C7",x"0019");
    gpmc_send('1',x"22C8",x"2700");
    gpmc_send('1',x"22C9",x"0018");
    gpmc_send('1',x"22CA",x"2800");
    gpmc_send('1',x"22CB",x"0017");
    gpmc_send('1',x"22CC",x"2900");
    gpmc_send('1',x"22CD",x"0016");
    gpmc_send('1',x"22CE",x"2A00");
    gpmc_send('1',x"22CF",x"0015");
    gpmc_send('1',x"22D0",x"2B00");
    gpmc_send('1',x"22D1",x"0014");
    gpmc_send('1',x"22D2",x"2C00");
    gpmc_send('1',x"22D3",x"0013");
    gpmc_send('1',x"22D4",x"2D00");
    gpmc_send('1',x"22D5",x"0012");
    gpmc_send('1',x"22D6",x"2E00");
    gpmc_send('1',x"22D7",x"0011");
    gpmc_send('1',x"22D8",x"2F00");
    gpmc_send('1',x"22D9",x"0010");
    gpmc_send('1',x"22DA",x"3000");
    gpmc_send('1',x"22DB",x"000F");
    gpmc_send('1',x"22DC",x"3100");
    gpmc_send('1',x"22DD",x"000E");
    gpmc_send('1',x"22DE",x"3200");
    gpmc_send('1',x"22DF",x"000D");
    gpmc_send('1',x"22E0",x"3300");
    gpmc_send('1',x"22E1",x"000C");
    gpmc_send('1',x"22E2",x"3400");
    gpmc_send('1',x"22E3",x"000B");
    gpmc_send('1',x"22E4",x"3500");
    gpmc_send('1',x"22E5",x"000A");
    gpmc_send('1',x"22E6",x"3600");
    gpmc_send('1',x"22E7",x"0009");
    gpmc_send('1',x"22E8",x"3700");
    gpmc_send('1',x"22E9",x"0008");
    gpmc_send('1',x"22EA",x"3800");
    gpmc_send('1',x"22EB",x"0007");
    gpmc_send('1',x"22EC",x"3900");
    gpmc_send('1',x"22ED",x"0006");
    gpmc_send('1',x"22EE",x"3A00");
    gpmc_send('1',x"22EF",x"0005");
    gpmc_send('1',x"22F0",x"3B00");
    gpmc_send('1',x"22F1",x"0004");
    gpmc_send('1',x"22F2",x"3C00");
    gpmc_send('1',x"22F3",x"0003");
    gpmc_send('1',x"22F4",x"3D00");
    gpmc_send('1',x"22F5",x"0002");
    gpmc_send('1',x"22F6",x"3E00");
    gpmc_send('1',x"22F7",x"0001");
    gpmc_send('1',x"22F8",x"3F00");
    gpmc_send('1',x"22F9",x"0000");
    gpmc_send('1',x"22FA",x"3F01");
    gpmc_send('1',x"22FB",x"0000");
    gpmc_send('1',x"22FC",x"3E02");
    gpmc_send('1',x"22FD",x"0000");
    gpmc_send('1',x"22FE",x"3D03");
    gpmc_send('1',x"22FF",x"0000");
    gpmc_send('1',x"2300",x"3C04");
    gpmc_send('1',x"2301",x"0000");
    gpmc_send('1',x"2302",x"3B05");
    gpmc_send('1',x"2303",x"0000");
    gpmc_send('1',x"2304",x"3A06");
    gpmc_send('1',x"2305",x"0000");
    gpmc_send('1',x"2306",x"3907");
    gpmc_send('1',x"2307",x"0000");
    gpmc_send('1',x"2308",x"3808");
    gpmc_send('1',x"2309",x"0000");
    gpmc_send('1',x"230A",x"3709");
    gpmc_send('1',x"230B",x"0000");
    gpmc_send('1',x"230C",x"360A");
    gpmc_send('1',x"230D",x"0000");
    gpmc_send('1',x"230E",x"350B");
    gpmc_send('1',x"230F",x"0000");
    gpmc_send('1',x"2310",x"340C");
    gpmc_send('1',x"2311",x"0000");
    gpmc_send('1',x"2312",x"330D");
    gpmc_send('1',x"2313",x"0000");
    gpmc_send('1',x"2314",x"320E");
    gpmc_send('1',x"2315",x"0000");
    gpmc_send('1',x"2316",x"310F");
    gpmc_send('1',x"2317",x"0000");
    gpmc_send('1',x"2318",x"3010");
    gpmc_send('1',x"2319",x"0000");
    gpmc_send('1',x"231A",x"2F11");
    gpmc_send('1',x"231B",x"0000");
    gpmc_send('1',x"231C",x"2E12");
    gpmc_send('1',x"231D",x"0000");
    gpmc_send('1',x"231E",x"2D13");
    gpmc_send('1',x"231F",x"0000");
    gpmc_send('1',x"2320",x"2C14");
    gpmc_send('1',x"2321",x"0000");
    gpmc_send('1',x"2322",x"2B15");
    gpmc_send('1',x"2323",x"0000");
    gpmc_send('1',x"2324",x"2A16");
    gpmc_send('1',x"2325",x"0000");
    gpmc_send('1',x"2326",x"2917");
    gpmc_send('1',x"2327",x"0000");
    gpmc_send('1',x"2328",x"2818");
    gpmc_send('1',x"2329",x"0000");
    gpmc_send('1',x"232A",x"2719");
    gpmc_send('1',x"232B",x"0000");
    gpmc_send('1',x"232C",x"261A");
    gpmc_send('1',x"232D",x"0000");
    gpmc_send('1',x"232E",x"251B");
    gpmc_send('1',x"232F",x"0000");
    gpmc_send('1',x"2330",x"241C");
    gpmc_send('1',x"2331",x"0000");
    gpmc_send('1',x"2332",x"231D");
    gpmc_send('1',x"2333",x"0000");
    gpmc_send('1',x"2334",x"221E");
    gpmc_send('1',x"2335",x"0000");
    gpmc_send('1',x"2336",x"211F");
    gpmc_send('1',x"2337",x"0000");
    gpmc_send('1',x"2338",x"2020");
    gpmc_send('1',x"2339",x"0000");
    gpmc_send('1',x"233A",x"1F21");
    gpmc_send('1',x"233B",x"0000");
    gpmc_send('1',x"233C",x"1E22");
    gpmc_send('1',x"233D",x"0000");
    gpmc_send('1',x"233E",x"1D23");
    gpmc_send('1',x"233F",x"0000");
    gpmc_send('1',x"2340",x"1C24");
    gpmc_send('1',x"2341",x"0000");
    gpmc_send('1',x"2342",x"1B25");
    gpmc_send('1',x"2343",x"0000");
    gpmc_send('1',x"2344",x"1A26");
    gpmc_send('1',x"2345",x"0000");
    gpmc_send('1',x"2346",x"1927");
    gpmc_send('1',x"2347",x"0000");
    gpmc_send('1',x"2348",x"1828");
    gpmc_send('1',x"2349",x"0000");
    gpmc_send('1',x"234A",x"1729");
    gpmc_send('1',x"234B",x"0000");
    gpmc_send('1',x"234C",x"162A");
    gpmc_send('1',x"234D",x"0000");
    gpmc_send('1',x"234E",x"152B");
    gpmc_send('1',x"234F",x"0000");
    gpmc_send('1',x"2350",x"142C");
    gpmc_send('1',x"2351",x"0000");
    gpmc_send('1',x"2352",x"132D");
    gpmc_send('1',x"2353",x"0000");
    gpmc_send('1',x"2354",x"122E");
    gpmc_send('1',x"2355",x"0000");
    gpmc_send('1',x"2356",x"112F");
    gpmc_send('1',x"2357",x"0000");
    gpmc_send('1',x"2358",x"1030");
    gpmc_send('1',x"2359",x"0000");
    gpmc_send('1',x"235A",x"0F31");
    gpmc_send('1',x"235B",x"0000");
    gpmc_send('1',x"235C",x"0E32");
    gpmc_send('1',x"235D",x"0000");
    gpmc_send('1',x"235E",x"0D33");
    gpmc_send('1',x"235F",x"0000");
    gpmc_send('1',x"2360",x"0C34");
    gpmc_send('1',x"2361",x"0000");
    gpmc_send('1',x"2362",x"0B35");
    gpmc_send('1',x"2363",x"0000");
    gpmc_send('1',x"2364",x"0A36");
    gpmc_send('1',x"2365",x"0000");
    gpmc_send('1',x"2366",x"0937");
    gpmc_send('1',x"2367",x"0000");
    gpmc_send('1',x"2368",x"0838");
    gpmc_send('1',x"2369",x"0000");
    gpmc_send('1',x"236A",x"0739");
    gpmc_send('1',x"236B",x"0000");
    gpmc_send('1',x"236C",x"063A");
    gpmc_send('1',x"236D",x"0000");
    gpmc_send('1',x"236E",x"053B");
    gpmc_send('1',x"236F",x"0000");
    gpmc_send('1',x"2370",x"043C");
    gpmc_send('1',x"2371",x"0000");
    gpmc_send('1',x"2372",x"033D");
    gpmc_send('1',x"2373",x"0000");
    gpmc_send('1',x"2374",x"023E");
    gpmc_send('1',x"2375",x"0000");
    gpmc_send('1',x"2376",x"013F");
    gpmc_send('1',x"2377",x"0000");
    gpmc_send('1',x"2378",x"003F");
    gpmc_send('1',x"2379",x"0000");
    gpmc_send('1',x"237A",x"003E");
    gpmc_send('1',x"237B",x"0001");
    gpmc_send('1',x"237C",x"003D");
    gpmc_send('1',x"237D",x"0002");
    gpmc_send('1',x"237E",x"003C");
    gpmc_send('1',x"237F",x"0003");
    gpmc_send('1',x"2380",x"003B");
    gpmc_send('1',x"2381",x"0004");
    gpmc_send('1',x"2382",x"003A");
    gpmc_send('1',x"2383",x"0005");
    gpmc_send('1',x"2384",x"0039");
    gpmc_send('1',x"2385",x"0006");
    gpmc_send('1',x"2386",x"0038");
    gpmc_send('1',x"2387",x"0007");
    gpmc_send('1',x"2388",x"0037");
    gpmc_send('1',x"2389",x"0008");
    gpmc_send('1',x"238A",x"0036");
    gpmc_send('1',x"238B",x"0009");
    gpmc_send('1',x"238C",x"0035");
    gpmc_send('1',x"238D",x"000A");
    gpmc_send('1',x"238E",x"0034");
    gpmc_send('1',x"238F",x"000B");
    gpmc_send('1',x"2390",x"0033");
    gpmc_send('1',x"2391",x"000C");
    gpmc_send('1',x"2392",x"0032");
    gpmc_send('1',x"2393",x"000D");
    gpmc_send('1',x"2394",x"0031");
    gpmc_send('1',x"2395",x"000E");
    gpmc_send('1',x"2396",x"0030");
    gpmc_send('1',x"2397",x"000F");
    gpmc_send('1',x"2398",x"002F");
    gpmc_send('1',x"2399",x"0010");
    gpmc_send('1',x"239A",x"002E");
    gpmc_send('1',x"239B",x"0011");
    gpmc_send('1',x"239C",x"002D");
    gpmc_send('1',x"239D",x"0012");
    gpmc_send('1',x"239E",x"002C");
    gpmc_send('1',x"239F",x"0013");
    gpmc_send('1',x"23A0",x"002B");
    gpmc_send('1',x"23A1",x"0014");
    gpmc_send('1',x"23A2",x"002A");
    gpmc_send('1',x"23A3",x"0015");
    gpmc_send('1',x"23A4",x"0029");
    gpmc_send('1',x"23A5",x"0016");
    gpmc_send('1',x"23A6",x"0028");
    gpmc_send('1',x"23A7",x"0017");
    gpmc_send('1',x"23A8",x"0027");
    gpmc_send('1',x"23A9",x"0018");
    gpmc_send('1',x"23AA",x"0026");
    gpmc_send('1',x"23AB",x"0019");
    gpmc_send('1',x"23AC",x"0025");
    gpmc_send('1',x"23AD",x"001A");
    gpmc_send('1',x"23AE",x"0024");
    gpmc_send('1',x"23AF",x"001B");
    gpmc_send('1',x"23B0",x"0023");
    gpmc_send('1',x"23B1",x"001C");
    gpmc_send('1',x"23B2",x"0022");
    gpmc_send('1',x"23B3",x"001D");
    gpmc_send('1',x"23B4",x"0021");
    gpmc_send('1',x"23B5",x"001E");
    gpmc_send('1',x"23B6",x"0020");
    gpmc_send('1',x"23B7",x"001F");
    gpmc_send('1',x"23B8",x"001F");
    gpmc_send('1',x"23B9",x"0020");
    gpmc_send('1',x"23BA",x"001E");
    gpmc_send('1',x"23BB",x"0021");
    gpmc_send('1',x"23BC",x"001D");
    gpmc_send('1',x"23BD",x"0022");
    gpmc_send('1',x"23BE",x"001C");
    gpmc_send('1',x"23BF",x"0023");
    gpmc_send('1',x"23C0",x"001B");
    gpmc_send('1',x"23C1",x"0024");
    gpmc_send('1',x"23C2",x"001A");
    gpmc_send('1',x"23C3",x"0025");
    gpmc_send('1',x"23C4",x"0019");
    gpmc_send('1',x"23C5",x"0026");
    gpmc_send('1',x"23C6",x"0018");
    gpmc_send('1',x"23C7",x"0027");
    gpmc_send('1',x"23C8",x"0017");
    gpmc_send('1',x"23C9",x"0028");
    gpmc_send('1',x"23CA",x"0016");
    gpmc_send('1',x"23CB",x"0029");
    gpmc_send('1',x"23CC",x"0015");
    gpmc_send('1',x"23CD",x"002A");
    gpmc_send('1',x"23CE",x"0014");
    gpmc_send('1',x"23CF",x"002B");
    gpmc_send('1',x"23D0",x"0013");
    gpmc_send('1',x"23D1",x"002C");
    gpmc_send('1',x"23D2",x"0012");
    gpmc_send('1',x"23D3",x"002D");
    gpmc_send('1',x"23D4",x"0011");
    gpmc_send('1',x"23D5",x"002E");
    gpmc_send('1',x"23D6",x"0010");
    gpmc_send('1',x"23D7",x"002F");
    gpmc_send('1',x"23D8",x"000F");
    gpmc_send('1',x"23D9",x"0030");
    gpmc_send('1',x"23DA",x"000E");
    gpmc_send('1',x"23DB",x"0031");
    gpmc_send('1',x"23DC",x"000D");
    gpmc_send('1',x"23DD",x"0032");
    gpmc_send('1',x"23DE",x"000C");
    gpmc_send('1',x"23DF",x"0033");
    gpmc_send('1',x"23E0",x"000B");
    gpmc_send('1',x"23E1",x"0034");
    gpmc_send('1',x"23E2",x"000A");
    gpmc_send('1',x"23E3",x"0035");
    gpmc_send('1',x"23E4",x"0009");
    gpmc_send('1',x"23E5",x"0036");
    gpmc_send('1',x"23E6",x"0008");
    gpmc_send('1',x"23E7",x"0037");
    gpmc_send('1',x"23E8",x"0007");
    gpmc_send('1',x"23E9",x"0038");
    gpmc_send('1',x"23EA",x"0006");
    gpmc_send('1',x"23EB",x"0039");
    gpmc_send('1',x"23EC",x"0005");
    gpmc_send('1',x"23ED",x"003A");
    gpmc_send('1',x"23EE",x"0004");
    gpmc_send('1',x"23EF",x"003B");
    gpmc_send('1',x"23F0",x"0003");
    gpmc_send('1',x"23F1",x"003C");
    gpmc_send('1',x"23F2",x"0002");
    gpmc_send('1',x"23F3",x"003D");
    gpmc_send('1',x"23F4",x"0001");
    gpmc_send('1',x"23F5",x"003E");
    gpmc_send('1',x"23F6",x"0000");
    gpmc_send('1',x"23F7",x"003F");
    gpmc_send('1',x"23F8",x"0100");
    gpmc_send('1',x"23F9",x"003E");
    gpmc_send('1',x"23FA",x"0200");
    gpmc_send('1',x"23FB",x"003D");
    gpmc_send('1',x"23FC",x"0300");
    gpmc_send('1',x"23FD",x"003C");
    gpmc_send('1',x"23FE",x"0400");
    gpmc_send('1',x"23FF",x"003B");
    gpmc_send('1',x"2400",x"0500");
    gpmc_send('1',x"2401",x"003A");
    gpmc_send('1',x"2402",x"0600");
    gpmc_send('1',x"2403",x"0039");
    gpmc_send('1',x"2404",x"0700");
    gpmc_send('1',x"2405",x"0038");
    gpmc_send('1',x"2406",x"0800");
    gpmc_send('1',x"2407",x"0037");
    gpmc_send('1',x"2408",x"0900");
    gpmc_send('1',x"2409",x"0036");
    gpmc_send('1',x"240A",x"0A00");
    gpmc_send('1',x"240B",x"0035");
    gpmc_send('1',x"240C",x"0B00");
    gpmc_send('1',x"240D",x"0034");
    gpmc_send('1',x"240E",x"0C00");
    gpmc_send('1',x"240F",x"0033");
    gpmc_send('1',x"2410",x"0D00");
    gpmc_send('1',x"2411",x"0032");
    gpmc_send('1',x"2412",x"0E00");
    gpmc_send('1',x"2413",x"0031");
    gpmc_send('1',x"2414",x"0F00");
    gpmc_send('1',x"2415",x"0030");
    gpmc_send('1',x"2416",x"1000");
    gpmc_send('1',x"2417",x"002F");
    gpmc_send('1',x"2418",x"1100");
    gpmc_send('1',x"2419",x"002E");
    gpmc_send('1',x"241A",x"1200");
    gpmc_send('1',x"241B",x"002D");
    gpmc_send('1',x"241C",x"1300");
    gpmc_send('1',x"241D",x"002C");
    gpmc_send('1',x"241E",x"1400");
    gpmc_send('1',x"241F",x"002B");
    gpmc_send('1',x"2420",x"1500");
    gpmc_send('1',x"2421",x"002A");
    gpmc_send('1',x"2422",x"1600");
    gpmc_send('1',x"2423",x"0029");
    gpmc_send('1',x"2424",x"1700");
    gpmc_send('1',x"2425",x"0028");
    gpmc_send('1',x"2426",x"1800");
    gpmc_send('1',x"2427",x"0027");
    gpmc_send('1',x"2428",x"1900");
    gpmc_send('1',x"2429",x"0026");
    gpmc_send('1',x"242A",x"1A00");
    gpmc_send('1',x"242B",x"0025");
    gpmc_send('1',x"242C",x"1B00");
    gpmc_send('1',x"242D",x"0024");
    gpmc_send('1',x"242E",x"1C00");
    gpmc_send('1',x"242F",x"0023");
    gpmc_send('1',x"2430",x"1D00");
    gpmc_send('1',x"2431",x"0022");
    gpmc_send('1',x"2432",x"1E00");
    gpmc_send('1',x"2433",x"0021");
    gpmc_send('1',x"2434",x"1F00");
    gpmc_send('1',x"2435",x"0020");
    gpmc_send('1',x"2436",x"2000");
    gpmc_send('1',x"2437",x"001F");
    gpmc_send('1',x"2438",x"2100");
    gpmc_send('1',x"2439",x"001E");
    gpmc_send('1',x"243A",x"2200");
    gpmc_send('1',x"243B",x"001D");
    gpmc_send('1',x"243C",x"2300");
    gpmc_send('1',x"243D",x"001C");
    gpmc_send('1',x"243E",x"2400");
    gpmc_send('1',x"243F",x"001B");
    gpmc_send('1',x"2440",x"2500");
    gpmc_send('1',x"2441",x"001A");
    gpmc_send('1',x"2442",x"2600");
    gpmc_send('1',x"2443",x"0019");
    gpmc_send('1',x"2444",x"2700");
    gpmc_send('1',x"2445",x"0018");
    gpmc_send('1',x"2446",x"2800");
    gpmc_send('1',x"2447",x"0017");
    gpmc_send('1',x"2448",x"2900");
    gpmc_send('1',x"2449",x"0016");
    gpmc_send('1',x"244A",x"2A00");
    gpmc_send('1',x"244B",x"0015");
    gpmc_send('1',x"244C",x"2B00");
    gpmc_send('1',x"244D",x"0014");
    gpmc_send('1',x"244E",x"2C00");
    gpmc_send('1',x"244F",x"0013");
    gpmc_send('1',x"2450",x"2D00");
    gpmc_send('1',x"2451",x"0012");
    gpmc_send('1',x"2452",x"2E00");
    gpmc_send('1',x"2453",x"0011");
    gpmc_send('1',x"2454",x"2F00");
    gpmc_send('1',x"2455",x"0010");
    gpmc_send('1',x"2456",x"3000");
    gpmc_send('1',x"2457",x"000F");
    gpmc_send('1',x"2458",x"3100");
    gpmc_send('1',x"2459",x"000E");
    gpmc_send('1',x"245A",x"3200");
    gpmc_send('1',x"245B",x"000D");
    gpmc_send('1',x"245C",x"3300");
    gpmc_send('1',x"245D",x"000C");
    gpmc_send('1',x"245E",x"3400");
    gpmc_send('1',x"245F",x"000B");
    gpmc_send('1',x"2460",x"3500");
    gpmc_send('1',x"2461",x"000A");
    gpmc_send('1',x"2462",x"3600");
    gpmc_send('1',x"2463",x"0009");
    gpmc_send('1',x"2464",x"3700");
    gpmc_send('1',x"2465",x"0008");
    gpmc_send('1',x"2466",x"3800");
    gpmc_send('1',x"2467",x"0007");
    gpmc_send('1',x"2468",x"3900");
    gpmc_send('1',x"2469",x"0006");
    gpmc_send('1',x"246A",x"3A00");
    gpmc_send('1',x"246B",x"0005");
    gpmc_send('1',x"246C",x"3B00");
    gpmc_send('1',x"246D",x"0004");
    gpmc_send('1',x"246E",x"3C00");
    gpmc_send('1',x"246F",x"0003");
    gpmc_send('1',x"2470",x"3D00");
    gpmc_send('1',x"2471",x"0002");
    gpmc_send('1',x"2472",x"3E00");
    gpmc_send('1',x"2473",x"0001");
    gpmc_send('1',x"2474",x"3F00");
    gpmc_send('1',x"2475",x"0000");
    gpmc_send('1',x"2476",x"3F01");
    gpmc_send('1',x"2477",x"0000");
    gpmc_send('1',x"2478",x"3E02");
    gpmc_send('1',x"2479",x"0000");
    gpmc_send('1',x"247A",x"3D03");
    gpmc_send('1',x"247B",x"0000");
    gpmc_send('1',x"247C",x"3C04");
    gpmc_send('1',x"247D",x"0000");
    gpmc_send('1',x"247E",x"3B05");
    gpmc_send('1',x"247F",x"0000");
    gpmc_send('1',x"2480",x"3A06");
    gpmc_send('1',x"2481",x"0000");
    gpmc_send('1',x"2482",x"3907");
    gpmc_send('1',x"2483",x"0000");
    gpmc_send('1',x"2484",x"3808");
    gpmc_send('1',x"2485",x"0000");
    gpmc_send('1',x"2486",x"3709");
    gpmc_send('1',x"2487",x"0000");
    gpmc_send('1',x"2488",x"360A");
    gpmc_send('1',x"2489",x"0000");
    gpmc_send('1',x"248A",x"350B");
    gpmc_send('1',x"248B",x"0000");
    gpmc_send('1',x"248C",x"340C");
    gpmc_send('1',x"248D",x"0000");
    gpmc_send('1',x"248E",x"330D");
    gpmc_send('1',x"248F",x"0000");
    gpmc_send('1',x"2490",x"320E");
    gpmc_send('1',x"2491",x"0000");
    gpmc_send('1',x"2492",x"310F");
    gpmc_send('1',x"2493",x"0000");
    gpmc_send('1',x"2494",x"3010");
    gpmc_send('1',x"2495",x"0000");
    gpmc_send('1',x"2496",x"2F11");
    gpmc_send('1',x"2497",x"0000");
    gpmc_send('1',x"2498",x"2E12");
    gpmc_send('1',x"2499",x"0000");
    gpmc_send('1',x"249A",x"2D13");
    gpmc_send('1',x"249B",x"0000");
    gpmc_send('1',x"249C",x"2C14");
    gpmc_send('1',x"249D",x"0000");
    gpmc_send('1',x"249E",x"2B15");
    gpmc_send('1',x"249F",x"0000");
    gpmc_send('1',x"24A0",x"2A16");
    gpmc_send('1',x"24A1",x"0000");
    gpmc_send('1',x"24A2",x"2917");
    gpmc_send('1',x"24A3",x"0000");
    gpmc_send('1',x"24A4",x"2818");
    gpmc_send('1',x"24A5",x"0000");
    gpmc_send('1',x"24A6",x"2719");
    gpmc_send('1',x"24A7",x"0000");
    gpmc_send('1',x"24A8",x"261A");
    gpmc_send('1',x"24A9",x"0000");
    gpmc_send('1',x"24AA",x"251B");
    gpmc_send('1',x"24AB",x"0000");
    gpmc_send('1',x"24AC",x"241C");
    gpmc_send('1',x"24AD",x"0000");
    gpmc_send('1',x"24AE",x"231D");
    gpmc_send('1',x"24AF",x"0000");
    gpmc_send('1',x"24B0",x"221E");
    gpmc_send('1',x"24B1",x"0000");
    gpmc_send('1',x"24B2",x"211F");
    gpmc_send('1',x"24B3",x"0000");
    gpmc_send('1',x"24B4",x"2020");
    gpmc_send('1',x"24B5",x"0000");
    gpmc_send('1',x"24B6",x"1F21");
    gpmc_send('1',x"24B7",x"0000");
    gpmc_send('1',x"24B8",x"1E22");
    gpmc_send('1',x"24B9",x"0000");
    gpmc_send('1',x"24BA",x"1D23");
    gpmc_send('1',x"24BB",x"0000");
    gpmc_send('1',x"24BC",x"1C24");
    gpmc_send('1',x"24BD",x"0000");
    gpmc_send('1',x"24BE",x"1B25");
    gpmc_send('1',x"24BF",x"0000");
    gpmc_send('1',x"24C0",x"1A26");
    gpmc_send('1',x"24C1",x"0000");
    gpmc_send('1',x"24C2",x"1927");
    gpmc_send('1',x"24C3",x"0000");
    gpmc_send('1',x"24C4",x"1828");
    gpmc_send('1',x"24C5",x"0000");
    gpmc_send('1',x"24C6",x"1729");
    gpmc_send('1',x"24C7",x"0000");
    gpmc_send('1',x"24C8",x"162A");
    gpmc_send('1',x"24C9",x"0000");
    gpmc_send('1',x"24CA",x"152B");
    gpmc_send('1',x"24CB",x"0000");
    gpmc_send('1',x"24CC",x"142C");
    gpmc_send('1',x"24CD",x"0000");
    gpmc_send('1',x"24CE",x"132D");
    gpmc_send('1',x"24CF",x"0000");
    gpmc_send('1',x"24D0",x"122E");
    gpmc_send('1',x"24D1",x"0000");
    gpmc_send('1',x"24D2",x"112F");
    gpmc_send('1',x"24D3",x"0000");
    gpmc_send('1',x"24D4",x"1030");
    gpmc_send('1',x"24D5",x"0000");
    gpmc_send('1',x"24D6",x"0F31");
    gpmc_send('1',x"24D7",x"0000");
    gpmc_send('1',x"24D8",x"0E32");
    gpmc_send('1',x"24D9",x"0000");
    gpmc_send('1',x"24DA",x"0D33");
    gpmc_send('1',x"24DB",x"0000");
    gpmc_send('1',x"24DC",x"0C34");
    gpmc_send('1',x"24DD",x"0000");
    gpmc_send('1',x"24DE",x"0B35");
    gpmc_send('1',x"24DF",x"0000");
    gpmc_send('1',x"24E0",x"0A36");
    gpmc_send('1',x"24E1",x"0000");
    gpmc_send('1',x"24E2",x"0937");
    gpmc_send('1',x"24E3",x"0000");
    gpmc_send('1',x"24E4",x"0838");
    gpmc_send('1',x"24E5",x"0000");
    gpmc_send('1',x"24E6",x"0739");
    gpmc_send('1',x"24E7",x"0000");
    gpmc_send('1',x"24E8",x"063A");
    gpmc_send('1',x"24E9",x"0000");
    gpmc_send('1',x"24EA",x"053B");
    gpmc_send('1',x"24EB",x"0000");
    gpmc_send('1',x"24EC",x"043C");
    gpmc_send('1',x"24ED",x"0000");
    gpmc_send('1',x"24EE",x"033D");
    gpmc_send('1',x"24EF",x"0000");
    gpmc_send('1',x"24F0",x"023E");
    gpmc_send('1',x"24F1",x"0000");
    gpmc_send('1',x"24F2",x"013F");
    gpmc_send('1',x"24F3",x"0000");
    gpmc_send('1',x"24F4",x"003F");
    gpmc_send('1',x"24F5",x"0000");
    gpmc_send('1',x"24F6",x"003E");
    gpmc_send('1',x"24F7",x"0001");
    gpmc_send('1',x"24F8",x"003D");
    gpmc_send('1',x"24F9",x"0002");
    gpmc_send('1',x"24FA",x"003C");
    gpmc_send('1',x"24FB",x"0003");
    gpmc_send('1',x"24FC",x"003B");
    gpmc_send('1',x"24FD",x"0004");
    gpmc_send('1',x"24FE",x"003A");
    gpmc_send('1',x"24FF",x"0005");
    gpmc_send('1',x"2500",x"0039");
    gpmc_send('1',x"2501",x"0006");
    gpmc_send('1',x"2502",x"0038");
    gpmc_send('1',x"2503",x"0007");
    gpmc_send('1',x"2504",x"0037");
    gpmc_send('1',x"2505",x"0008");
    gpmc_send('1',x"2506",x"0036");
    gpmc_send('1',x"2507",x"0009");
    gpmc_send('1',x"2508",x"0035");
    gpmc_send('1',x"2509",x"000A");
    gpmc_send('1',x"250A",x"0034");
    gpmc_send('1',x"250B",x"000B");
    gpmc_send('1',x"250C",x"0033");
    gpmc_send('1',x"250D",x"000C");
    gpmc_send('1',x"250E",x"0032");
    gpmc_send('1',x"250F",x"000D");
    gpmc_send('1',x"2510",x"0031");
    gpmc_send('1',x"2511",x"000E");
    gpmc_send('1',x"2512",x"0030");
    gpmc_send('1',x"2513",x"000F");
    gpmc_send('1',x"2514",x"002F");
    gpmc_send('1',x"2515",x"0010");
    gpmc_send('1',x"2516",x"002E");
    gpmc_send('1',x"2517",x"0011");
    gpmc_send('1',x"2518",x"002D");
    gpmc_send('1',x"2519",x"0012");
    gpmc_send('1',x"251A",x"002C");
    gpmc_send('1',x"251B",x"0013");
    gpmc_send('1',x"251C",x"002B");
    gpmc_send('1',x"251D",x"0014");
    gpmc_send('1',x"251E",x"002A");
    gpmc_send('1',x"251F",x"0015");
    gpmc_send('1',x"2520",x"0029");
    gpmc_send('1',x"2521",x"0016");
    gpmc_send('1',x"2522",x"0028");
    gpmc_send('1',x"2523",x"0017");
    gpmc_send('1',x"2524",x"0027");
    gpmc_send('1',x"2525",x"0018");
    gpmc_send('1',x"2526",x"0026");
    gpmc_send('1',x"2527",x"0019");
    gpmc_send('1',x"2528",x"0025");
    gpmc_send('1',x"2529",x"001A");
    gpmc_send('1',x"252A",x"0024");
    gpmc_send('1',x"252B",x"001B");
    gpmc_send('1',x"252C",x"0023");
    gpmc_send('1',x"252D",x"001C");
    gpmc_send('1',x"252E",x"0022");
    gpmc_send('1',x"252F",x"001D");
    gpmc_send('1',x"2530",x"0021");
    gpmc_send('1',x"2531",x"001E");
    gpmc_send('1',x"2532",x"0020");
    gpmc_send('1',x"2533",x"001F");
    gpmc_send('1',x"2534",x"001F");
    gpmc_send('1',x"2535",x"0020");
    gpmc_send('1',x"2536",x"001E");
    gpmc_send('1',x"2537",x"0021");
    gpmc_send('1',x"2538",x"001D");
    gpmc_send('1',x"2539",x"0022");
    gpmc_send('1',x"253A",x"001C");
    gpmc_send('1',x"253B",x"0023");
    gpmc_send('1',x"253C",x"001B");
    gpmc_send('1',x"253D",x"0024");
    gpmc_send('1',x"253E",x"001A");
    gpmc_send('1',x"253F",x"0025");
    gpmc_send('1',x"2540",x"0019");
    gpmc_send('1',x"2541",x"0026");
    gpmc_send('1',x"2542",x"0018");
    gpmc_send('1',x"2543",x"0027");
    gpmc_send('1',x"2544",x"0017");
    gpmc_send('1',x"2545",x"0028");
    gpmc_send('1',x"2546",x"0016");
    gpmc_send('1',x"2547",x"0029");
    gpmc_send('1',x"2548",x"0015");
    gpmc_send('1',x"2549",x"002A");
    gpmc_send('1',x"254A",x"0014");
    gpmc_send('1',x"254B",x"002B");
    gpmc_send('1',x"254C",x"0013");
    gpmc_send('1',x"254D",x"002C");
    gpmc_send('1',x"254E",x"0012");
    gpmc_send('1',x"254F",x"002D");
    gpmc_send('1',x"2550",x"0011");
    gpmc_send('1',x"2551",x"002E");
    gpmc_send('1',x"2552",x"0010");
    gpmc_send('1',x"2553",x"002F");
    gpmc_send('1',x"2554",x"000F");
    gpmc_send('1',x"2555",x"0030");
    gpmc_send('1',x"2556",x"000E");
    gpmc_send('1',x"2557",x"0031");
    gpmc_send('1',x"2558",x"000D");
    gpmc_send('1',x"2559",x"0032");
    gpmc_send('1',x"255A",x"000C");
    gpmc_send('1',x"255B",x"0033");
    gpmc_send('1',x"255C",x"000B");
    gpmc_send('1',x"255D",x"0034");
    gpmc_send('1',x"255E",x"000A");
    gpmc_send('1',x"255F",x"0035");
    gpmc_send('1',x"2560",x"0009");
    gpmc_send('1',x"2561",x"0036");
    gpmc_send('1',x"2562",x"0008");
    gpmc_send('1',x"2563",x"0037");
    gpmc_send('1',x"2564",x"0007");
    gpmc_send('1',x"2565",x"0038");
    gpmc_send('1',x"2566",x"0006");
    gpmc_send('1',x"2567",x"0039");
    gpmc_send('1',x"2568",x"0005");
    gpmc_send('1',x"2569",x"003A");
    gpmc_send('1',x"256A",x"0004");
    gpmc_send('1',x"256B",x"003B");
    gpmc_send('1',x"256C",x"0003");
    gpmc_send('1',x"256D",x"003C");
    gpmc_send('1',x"256E",x"0002");
    gpmc_send('1',x"256F",x"003D");
    gpmc_send('1',x"2570",x"0001");
    gpmc_send('1',x"2571",x"003E");
    gpmc_send('1',x"2572",x"0000");
    gpmc_send('1',x"2573",x"003F");
    gpmc_send('1',x"2574",x"0100");
    gpmc_send('1',x"2575",x"003E");
    gpmc_send('1',x"2576",x"0200");
    gpmc_send('1',x"2577",x"003D");
    gpmc_send('1',x"2578",x"0300");
    gpmc_send('1',x"2579",x"003C");
    gpmc_send('1',x"257A",x"0400");
    gpmc_send('1',x"257B",x"003B");
    gpmc_send('1',x"257C",x"0500");
    gpmc_send('1',x"257D",x"003A");
    gpmc_send('1',x"257E",x"0600");
    gpmc_send('1',x"257F",x"0039");
    gpmc_send('1',x"2580",x"0700");
    gpmc_send('1',x"2581",x"0038");
    gpmc_send('1',x"2582",x"0800");
    gpmc_send('1',x"2583",x"0037");
    gpmc_send('1',x"2584",x"0900");
    gpmc_send('1',x"2585",x"0036");
    gpmc_send('1',x"2586",x"0A00");
    gpmc_send('1',x"2587",x"0035");
    gpmc_send('1',x"2588",x"0B00");
    gpmc_send('1',x"2589",x"0034");
    gpmc_send('1',x"258A",x"0C00");
    gpmc_send('1',x"258B",x"0033");
    gpmc_send('1',x"258C",x"0D00");
    gpmc_send('1',x"258D",x"0032");
    gpmc_send('1',x"258E",x"0E00");
    gpmc_send('1',x"258F",x"0031");
    gpmc_send('1',x"2590",x"0F00");
    gpmc_send('1',x"2591",x"0030");
    gpmc_send('1',x"2592",x"1000");
    gpmc_send('1',x"2593",x"002F");
    gpmc_send('1',x"2594",x"1100");
    gpmc_send('1',x"2595",x"002E");
    gpmc_send('1',x"2596",x"1200");
    gpmc_send('1',x"2597",x"002D");
    gpmc_send('1',x"2598",x"1300");
    gpmc_send('1',x"2599",x"002C");
    gpmc_send('1',x"259A",x"1400");
    gpmc_send('1',x"259B",x"002B");
    gpmc_send('1',x"259C",x"1500");
    gpmc_send('1',x"259D",x"002A");
    gpmc_send('1',x"259E",x"1600");
    gpmc_send('1',x"259F",x"0029");
    gpmc_send('1',x"25A0",x"1700");
    gpmc_send('1',x"25A1",x"0028");
    gpmc_send('1',x"25A2",x"1800");
    gpmc_send('1',x"25A3",x"0027");
    gpmc_send('1',x"25A4",x"1900");
    gpmc_send('1',x"25A5",x"0026");
    gpmc_send('1',x"25A6",x"1A00");
    gpmc_send('1',x"25A7",x"0025");
    gpmc_send('1',x"25A8",x"1B00");
    gpmc_send('1',x"25A9",x"0024");
    gpmc_send('1',x"25AA",x"1C00");
    gpmc_send('1',x"25AB",x"0023");
    gpmc_send('1',x"25AC",x"1D00");
    gpmc_send('1',x"25AD",x"0022");
    gpmc_send('1',x"25AE",x"1E00");
    gpmc_send('1',x"25AF",x"0021");
    gpmc_send('1',x"25B0",x"1F00");
    gpmc_send('1',x"25B1",x"0020");
    gpmc_send('1',x"25B2",x"2000");
    gpmc_send('1',x"25B3",x"001F");
    gpmc_send('1',x"25B4",x"2100");
    gpmc_send('1',x"25B5",x"001E");
    gpmc_send('1',x"25B6",x"2200");
    gpmc_send('1',x"25B7",x"001D");
    gpmc_send('1',x"25B8",x"2300");
    gpmc_send('1',x"25B9",x"001C");
    gpmc_send('1',x"25BA",x"2400");
    gpmc_send('1',x"25BB",x"001B");
    gpmc_send('1',x"25BC",x"2500");
    gpmc_send('1',x"25BD",x"001A");
    gpmc_send('1',x"25BE",x"2600");
    gpmc_send('1',x"25BF",x"0019");
    gpmc_send('1',x"25C0",x"2700");
    gpmc_send('1',x"25C1",x"0018");
    gpmc_send('1',x"25C2",x"2800");
    gpmc_send('1',x"25C3",x"0017");
    gpmc_send('1',x"25C4",x"2900");
    gpmc_send('1',x"25C5",x"0016");
    gpmc_send('1',x"25C6",x"2A00");
    gpmc_send('1',x"25C7",x"0015");
    gpmc_send('1',x"25C8",x"2B00");
    gpmc_send('1',x"25C9",x"0014");
    gpmc_send('1',x"25CA",x"2C00");
    gpmc_send('1',x"25CB",x"0013");
    gpmc_send('1',x"25CC",x"2D00");
    gpmc_send('1',x"25CD",x"0012");
    gpmc_send('1',x"25CE",x"2E00");
    gpmc_send('1',x"25CF",x"0011");
    gpmc_send('1',x"25D0",x"2F00");
    gpmc_send('1',x"25D1",x"0010");
    gpmc_send('1',x"25D2",x"3000");
    gpmc_send('1',x"25D3",x"000F");
    gpmc_send('1',x"25D4",x"3100");
    gpmc_send('1',x"25D5",x"000E");
    gpmc_send('1',x"25D6",x"3200");
    gpmc_send('1',x"25D7",x"000D");
    gpmc_send('1',x"25D8",x"3300");
    gpmc_send('1',x"25D9",x"000C");
    gpmc_send('1',x"25DA",x"3400");
    gpmc_send('1',x"25DB",x"000B");
    gpmc_send('1',x"25DC",x"3500");
    gpmc_send('1',x"25DD",x"000A");
    gpmc_send('1',x"25DE",x"3600");
    gpmc_send('1',x"25DF",x"0009");
    gpmc_send('1',x"25E0",x"3700");
    gpmc_send('1',x"25E1",x"0008");
    gpmc_send('1',x"25E2",x"3800");
    gpmc_send('1',x"25E3",x"0007");
    gpmc_send('1',x"25E4",x"3900");
    gpmc_send('1',x"25E5",x"0006");
    gpmc_send('1',x"25E6",x"3A00");
    gpmc_send('1',x"25E7",x"0005");
    gpmc_send('1',x"25E8",x"3B00");
    gpmc_send('1',x"25E9",x"0004");
    gpmc_send('1',x"25EA",x"3C00");
    gpmc_send('1',x"25EB",x"0003");
    gpmc_send('1',x"25EC",x"3D00");
    gpmc_send('1',x"25ED",x"0002");
    gpmc_send('1',x"25EE",x"3E00");
    gpmc_send('1',x"25EF",x"0001");
    gpmc_send('1',x"25F0",x"3F00");
    gpmc_send('1',x"25F1",x"0000");
    gpmc_send('1',x"25F2",x"3F01");
    gpmc_send('1',x"25F3",x"0000");
    gpmc_send('1',x"25F4",x"3E02");
    gpmc_send('1',x"25F5",x"0000");
    gpmc_send('1',x"25F6",x"3D03");
    gpmc_send('1',x"25F7",x"0000");
    gpmc_send('1',x"25F8",x"3C04");
    gpmc_send('1',x"25F9",x"0000");
    gpmc_send('1',x"25FA",x"3B05");
    gpmc_send('1',x"25FB",x"0000");
    gpmc_send('1',x"25FC",x"3A06");
    gpmc_send('1',x"25FD",x"0000");
    gpmc_send('1',x"25FE",x"3907");
    gpmc_send('1',x"25FF",x"0000");
    gpmc_send('1',x"2600",x"3808");
    gpmc_send('1',x"2601",x"0000");
    gpmc_send('1',x"2602",x"3709");
    gpmc_send('1',x"2603",x"0000");
    gpmc_send('1',x"2604",x"360A");
    gpmc_send('1',x"2605",x"0000");
    gpmc_send('1',x"2606",x"350B");
    gpmc_send('1',x"2607",x"0000");
    gpmc_send('1',x"2608",x"340C");
    gpmc_send('1',x"2609",x"0000");
    gpmc_send('1',x"260A",x"330D");
    gpmc_send('1',x"260B",x"0000");
    gpmc_send('1',x"260C",x"320E");
    gpmc_send('1',x"260D",x"0000");
    gpmc_send('1',x"260E",x"310F");
    gpmc_send('1',x"260F",x"0000");
    gpmc_send('1',x"2610",x"3010");
    gpmc_send('1',x"2611",x"0000");
    gpmc_send('1',x"2612",x"2F11");
    gpmc_send('1',x"2613",x"0000");
    gpmc_send('1',x"2614",x"2E12");
    gpmc_send('1',x"2615",x"0000");
    gpmc_send('1',x"2616",x"2D13");
    gpmc_send('1',x"2617",x"0000");
    gpmc_send('1',x"2618",x"2C14");
    gpmc_send('1',x"2619",x"0000");
    gpmc_send('1',x"261A",x"2B15");
    gpmc_send('1',x"261B",x"0000");
    gpmc_send('1',x"261C",x"2A16");
    gpmc_send('1',x"261D",x"0000");
    gpmc_send('1',x"261E",x"2917");
    gpmc_send('1',x"261F",x"0000");
    gpmc_send('1',x"2620",x"2818");
    gpmc_send('1',x"2621",x"0000");
    gpmc_send('1',x"2622",x"2719");
    gpmc_send('1',x"2623",x"0000");
    gpmc_send('1',x"2624",x"261A");
    gpmc_send('1',x"2625",x"0000");
    gpmc_send('1',x"2626",x"251B");
    gpmc_send('1',x"2627",x"0000");
    gpmc_send('1',x"2628",x"241C");
    gpmc_send('1',x"2629",x"0000");
    gpmc_send('1',x"262A",x"231D");
    gpmc_send('1',x"262B",x"0000");
    gpmc_send('1',x"262C",x"221E");
    gpmc_send('1',x"262D",x"0000");
    gpmc_send('1',x"262E",x"211F");
    gpmc_send('1',x"262F",x"0000");
    gpmc_send('1',x"2630",x"2020");
    gpmc_send('1',x"2631",x"0000");
    gpmc_send('1',x"2632",x"1F21");
    gpmc_send('1',x"2633",x"0000");
    gpmc_send('1',x"2634",x"1E22");
    gpmc_send('1',x"2635",x"0000");
    gpmc_send('1',x"2636",x"1D23");
    gpmc_send('1',x"2637",x"0000");
    gpmc_send('1',x"2638",x"1C24");
    gpmc_send('1',x"2639",x"0000");
    gpmc_send('1',x"263A",x"1B25");
    gpmc_send('1',x"263B",x"0000");
    gpmc_send('1',x"263C",x"1A26");
    gpmc_send('1',x"263D",x"0000");
    gpmc_send('1',x"263E",x"1927");
    gpmc_send('1',x"263F",x"0000");
    gpmc_send('1',x"2640",x"1828");
    gpmc_send('1',x"2641",x"0000");
    gpmc_send('1',x"2642",x"1729");
    gpmc_send('1',x"2643",x"0000");
    gpmc_send('1',x"2644",x"162A");
    gpmc_send('1',x"2645",x"0000");
    gpmc_send('1',x"2646",x"152B");
    gpmc_send('1',x"2647",x"0000");
    gpmc_send('1',x"2648",x"142C");
    gpmc_send('1',x"2649",x"0000");
    gpmc_send('1',x"264A",x"132D");
    gpmc_send('1',x"264B",x"0000");
    gpmc_send('1',x"264C",x"122E");
    gpmc_send('1',x"264D",x"0000");
    gpmc_send('1',x"264E",x"112F");
    gpmc_send('1',x"264F",x"0000");
    gpmc_send('1',x"2650",x"1030");
    gpmc_send('1',x"2651",x"0000");
    gpmc_send('1',x"2652",x"0F31");
    gpmc_send('1',x"2653",x"0000");
    gpmc_send('1',x"2654",x"0E32");
    gpmc_send('1',x"2655",x"0000");
    gpmc_send('1',x"2656",x"0D33");
    gpmc_send('1',x"2657",x"0000");
    gpmc_send('1',x"2658",x"0C34");
    gpmc_send('1',x"2659",x"0000");
    gpmc_send('1',x"265A",x"0B35");
    gpmc_send('1',x"265B",x"0000");
    gpmc_send('1',x"265C",x"0A36");
    gpmc_send('1',x"265D",x"0000");
    gpmc_send('1',x"265E",x"0937");
    gpmc_send('1',x"265F",x"0000");
    gpmc_send('1',x"2660",x"0838");
    gpmc_send('1',x"2661",x"0000");
    gpmc_send('1',x"2662",x"0739");
    gpmc_send('1',x"2663",x"0000");
    gpmc_send('1',x"2664",x"063A");
    gpmc_send('1',x"2665",x"0000");
    gpmc_send('1',x"2666",x"053B");
    gpmc_send('1',x"2667",x"0000");
    gpmc_send('1',x"2668",x"043C");
    gpmc_send('1',x"2669",x"0000");
    gpmc_send('1',x"266A",x"033D");
    gpmc_send('1',x"266B",x"0000");
    gpmc_send('1',x"266C",x"023E");
    gpmc_send('1',x"266D",x"0000");
    gpmc_send('1',x"266E",x"013F");
    gpmc_send('1',x"266F",x"0000");
    gpmc_send('1',x"2670",x"003F");
    gpmc_send('1',x"2671",x"0000");
    gpmc_send('1',x"2672",x"003E");
    gpmc_send('1',x"2673",x"0001");
    gpmc_send('1',x"2674",x"003D");
    gpmc_send('1',x"2675",x"0002");
    gpmc_send('1',x"2676",x"003C");
    gpmc_send('1',x"2677",x"0003");
    gpmc_send('1',x"2678",x"003B");
    gpmc_send('1',x"2679",x"0004");
    gpmc_send('1',x"267A",x"003A");
    gpmc_send('1',x"267B",x"0005");
    gpmc_send('1',x"267C",x"0039");
    gpmc_send('1',x"267D",x"0006");
    gpmc_send('1',x"267E",x"0038");
    gpmc_send('1',x"267F",x"0007");
    gpmc_send('1',x"2680",x"0037");
    gpmc_send('1',x"2681",x"0008");
    gpmc_send('1',x"2682",x"0036");
    gpmc_send('1',x"2683",x"0009");
    gpmc_send('1',x"2684",x"0035");
    gpmc_send('1',x"2685",x"000A");
    gpmc_send('1',x"2686",x"0034");
    gpmc_send('1',x"2687",x"000B");
    gpmc_send('1',x"2688",x"0033");
    gpmc_send('1',x"2689",x"000C");
    gpmc_send('1',x"268A",x"0032");
    gpmc_send('1',x"268B",x"000D");
    gpmc_send('1',x"268C",x"0031");
    gpmc_send('1',x"268D",x"000E");
    gpmc_send('1',x"268E",x"0030");
    gpmc_send('1',x"268F",x"000F");
    gpmc_send('1',x"2690",x"002F");
    gpmc_send('1',x"2691",x"0010");
    gpmc_send('1',x"2692",x"002E");
    gpmc_send('1',x"2693",x"0011");
    gpmc_send('1',x"2694",x"002D");
    gpmc_send('1',x"2695",x"0012");
    gpmc_send('1',x"2696",x"002C");
    gpmc_send('1',x"2697",x"0013");
    gpmc_send('1',x"2698",x"002B");
    gpmc_send('1',x"2699",x"0014");
    gpmc_send('1',x"269A",x"002A");
    gpmc_send('1',x"269B",x"0015");
    gpmc_send('1',x"269C",x"0029");
    gpmc_send('1',x"269D",x"0016");
    gpmc_send('1',x"269E",x"0028");
    gpmc_send('1',x"269F",x"0017");
    gpmc_send('1',x"26A0",x"0027");
    gpmc_send('1',x"26A1",x"0018");
    gpmc_send('1',x"26A2",x"0026");
    gpmc_send('1',x"26A3",x"0019");
    gpmc_send('1',x"26A4",x"0025");
    gpmc_send('1',x"26A5",x"001A");
    gpmc_send('1',x"26A6",x"0024");
    gpmc_send('1',x"26A7",x"001B");
    gpmc_send('1',x"26A8",x"0023");
    gpmc_send('1',x"26A9",x"001C");
    gpmc_send('1',x"26AA",x"0022");
    gpmc_send('1',x"26AB",x"001D");
    gpmc_send('1',x"26AC",x"0021");
    gpmc_send('1',x"26AD",x"001E");
    gpmc_send('1',x"26AE",x"0020");
    gpmc_send('1',x"26AF",x"001F");
    gpmc_send('1',x"26B0",x"001F");
    gpmc_send('1',x"26B1",x"0020");
    gpmc_send('1',x"26B2",x"001E");
    gpmc_send('1',x"26B3",x"0021");
    gpmc_send('1',x"26B4",x"001D");
    gpmc_send('1',x"26B5",x"0022");
    gpmc_send('1',x"26B6",x"001C");
    gpmc_send('1',x"26B7",x"0023");
    gpmc_send('1',x"26B8",x"001B");
    gpmc_send('1',x"26B9",x"0024");
    gpmc_send('1',x"26BA",x"001A");
    gpmc_send('1',x"26BB",x"0025");
    gpmc_send('1',x"26BC",x"0019");
    gpmc_send('1',x"26BD",x"0026");
    gpmc_send('1',x"26BE",x"0018");
    gpmc_send('1',x"26BF",x"0027");
    gpmc_send('1',x"26C0",x"0017");
    gpmc_send('1',x"26C1",x"0028");
    gpmc_send('1',x"26C2",x"0016");
    gpmc_send('1',x"26C3",x"0029");
    gpmc_send('1',x"26C4",x"0015");
    gpmc_send('1',x"26C5",x"002A");
    gpmc_send('1',x"26C6",x"0014");
    gpmc_send('1',x"26C7",x"002B");
    gpmc_send('1',x"26C8",x"0013");
    gpmc_send('1',x"26C9",x"002C");
    gpmc_send('1',x"26CA",x"0012");
    gpmc_send('1',x"26CB",x"002D");
    gpmc_send('1',x"26CC",x"0011");
    gpmc_send('1',x"26CD",x"002E");
    gpmc_send('1',x"26CE",x"0010");
    gpmc_send('1',x"26CF",x"002F");
    gpmc_send('1',x"26D0",x"000F");
    gpmc_send('1',x"26D1",x"0030");
    gpmc_send('1',x"26D2",x"000E");
    gpmc_send('1',x"26D3",x"0031");
    gpmc_send('1',x"26D4",x"000D");
    gpmc_send('1',x"26D5",x"0032");
    gpmc_send('1',x"26D6",x"000C");
    gpmc_send('1',x"26D7",x"0033");
    gpmc_send('1',x"26D8",x"000B");
    gpmc_send('1',x"26D9",x"0034");
    gpmc_send('1',x"26DA",x"000A");
    gpmc_send('1',x"26DB",x"0035");
    gpmc_send('1',x"26DC",x"0009");
    gpmc_send('1',x"26DD",x"0036");
    gpmc_send('1',x"26DE",x"0008");
    gpmc_send('1',x"26DF",x"0037");
    gpmc_send('1',x"26E0",x"0007");
    gpmc_send('1',x"26E1",x"0038");
    gpmc_send('1',x"26E2",x"0006");
    gpmc_send('1',x"26E3",x"0039");
    gpmc_send('1',x"26E4",x"0005");
    gpmc_send('1',x"26E5",x"003A");
    gpmc_send('1',x"26E6",x"0004");
    gpmc_send('1',x"26E7",x"003B");
    gpmc_send('1',x"26E8",x"0003");
    gpmc_send('1',x"26E9",x"003C");
    gpmc_send('1',x"26EA",x"0002");
    gpmc_send('1',x"26EB",x"003D");
    gpmc_send('1',x"26EC",x"0001");
    gpmc_send('1',x"26ED",x"003E");
    gpmc_send('1',x"26EE",x"0000");
    gpmc_send('1',x"26EF",x"003F");
    gpmc_send('1',x"26F0",x"0100");
    gpmc_send('1',x"26F1",x"003E");
    gpmc_send('1',x"26F2",x"0200");
    gpmc_send('1',x"26F3",x"003D");
    gpmc_send('1',x"26F4",x"0300");
    gpmc_send('1',x"26F5",x"003C");
    gpmc_send('1',x"26F6",x"0400");
    gpmc_send('1',x"26F7",x"003B");
    gpmc_send('1',x"26F8",x"0500");
    gpmc_send('1',x"26F9",x"003A");
    gpmc_send('1',x"26FA",x"0600");
    gpmc_send('1',x"26FB",x"0039");
    gpmc_send('1',x"26FC",x"0700");
    gpmc_send('1',x"26FD",x"0038");
    gpmc_send('1',x"26FE",x"0800");
    gpmc_send('1',x"26FF",x"0037");
    gpmc_send('1',x"2700",x"0900");
    gpmc_send('1',x"2701",x"0036");
    gpmc_send('1',x"2702",x"0A00");
    gpmc_send('1',x"2703",x"0035");
    gpmc_send('1',x"2704",x"0B00");
    gpmc_send('1',x"2705",x"0034");
    gpmc_send('1',x"2706",x"0C00");
    gpmc_send('1',x"2707",x"0033");
    gpmc_send('1',x"2708",x"0D00");
    gpmc_send('1',x"2709",x"0032");
    gpmc_send('1',x"270A",x"0E00");
    gpmc_send('1',x"270B",x"0031");
    gpmc_send('1',x"270C",x"0F00");
    gpmc_send('1',x"270D",x"0030");
    gpmc_send('1',x"270E",x"1000");
    gpmc_send('1',x"270F",x"002F");
    gpmc_send('1',x"2710",x"1100");
    gpmc_send('1',x"2711",x"002E");
    gpmc_send('1',x"2712",x"1200");
    gpmc_send('1',x"2713",x"002D");
    gpmc_send('1',x"2714",x"1300");
    gpmc_send('1',x"2715",x"002C");
    gpmc_send('1',x"2716",x"1400");
    gpmc_send('1',x"2717",x"002B");
    gpmc_send('1',x"2718",x"1500");
    gpmc_send('1',x"2719",x"002A");
    gpmc_send('1',x"271A",x"1600");
    gpmc_send('1',x"271B",x"0029");
    gpmc_send('1',x"271C",x"1700");
    gpmc_send('1',x"271D",x"0028");
    gpmc_send('1',x"271E",x"1800");
    gpmc_send('1',x"271F",x"0027");
    gpmc_send('1',x"2720",x"1900");
    gpmc_send('1',x"2721",x"0026");
    gpmc_send('1',x"2722",x"1A00");
    gpmc_send('1',x"2723",x"0025");
    gpmc_send('1',x"2724",x"1B00");
    gpmc_send('1',x"2725",x"0024");
    gpmc_send('1',x"2726",x"1C00");
    gpmc_send('1',x"2727",x"0023");
    gpmc_send('1',x"2728",x"1D00");
    gpmc_send('1',x"2729",x"0022");
    gpmc_send('1',x"272A",x"1E00");
    gpmc_send('1',x"272B",x"0021");
    gpmc_send('1',x"272C",x"1F00");
    gpmc_send('1',x"272D",x"0020");
    gpmc_send('1',x"272E",x"2000");
    gpmc_send('1',x"272F",x"001F");
    gpmc_send('1',x"2730",x"2100");
    gpmc_send('1',x"2731",x"001E");
    gpmc_send('1',x"2732",x"2200");
    gpmc_send('1',x"2733",x"001D");
    gpmc_send('1',x"2734",x"2300");
    gpmc_send('1',x"2735",x"001C");
    gpmc_send('1',x"2736",x"2400");
    gpmc_send('1',x"2737",x"001B");
    gpmc_send('1',x"2738",x"2500");
    gpmc_send('1',x"2739",x"001A");
    gpmc_send('1',x"273A",x"2600");
    gpmc_send('1',x"273B",x"0019");
    gpmc_send('1',x"273C",x"2700");
    gpmc_send('1',x"273D",x"0018");
    gpmc_send('1',x"273E",x"2800");
    gpmc_send('1',x"273F",x"0017");
    gpmc_send('1',x"2740",x"2900");
    gpmc_send('1',x"2741",x"0016");
    gpmc_send('1',x"2742",x"2A00");
    gpmc_send('1',x"2743",x"0015");
    gpmc_send('1',x"2744",x"2B00");
    gpmc_send('1',x"2745",x"0014");
    gpmc_send('1',x"2746",x"2C00");
    gpmc_send('1',x"2747",x"0013");
    gpmc_send('1',x"2748",x"2D00");
    gpmc_send('1',x"2749",x"0012");
    gpmc_send('1',x"274A",x"2E00");
    gpmc_send('1',x"274B",x"0011");
    gpmc_send('1',x"274C",x"2F00");
    gpmc_send('1',x"274D",x"0010");
    gpmc_send('1',x"274E",x"3000");
    gpmc_send('1',x"274F",x"000F");
    gpmc_send('1',x"2750",x"3100");
    gpmc_send('1',x"2751",x"000E");
    gpmc_send('1',x"2752",x"3200");
    gpmc_send('1',x"2753",x"000D");
    gpmc_send('1',x"2754",x"3300");
    gpmc_send('1',x"2755",x"000C");
    gpmc_send('1',x"2756",x"3400");
    gpmc_send('1',x"2757",x"000B");
    gpmc_send('1',x"2758",x"3500");
    gpmc_send('1',x"2759",x"000A");
    gpmc_send('1',x"275A",x"3600");
    gpmc_send('1',x"275B",x"0009");
    gpmc_send('1',x"275C",x"3700");
    gpmc_send('1',x"275D",x"0008");
    gpmc_send('1',x"275E",x"3800");
    gpmc_send('1',x"275F",x"0007");
    gpmc_send('1',x"2760",x"3900");
    gpmc_send('1',x"2761",x"0006");
    gpmc_send('1',x"2762",x"3A00");
    gpmc_send('1',x"2763",x"0005");
    gpmc_send('1',x"2764",x"3B00");
    gpmc_send('1',x"2765",x"0004");
    gpmc_send('1',x"2766",x"3C00");
    gpmc_send('1',x"2767",x"0003");
    gpmc_send('1',x"2768",x"3D00");
    gpmc_send('1',x"2769",x"0002");
    gpmc_send('1',x"276A",x"3E00");
    gpmc_send('1',x"276B",x"0001");
    gpmc_send('1',x"276C",x"3F00");
    gpmc_send('1',x"276D",x"0000");
    gpmc_send('1',x"276E",x"3F01");
    gpmc_send('1',x"276F",x"0000");
    gpmc_send('1',x"2770",x"3E02");
    gpmc_send('1',x"2771",x"0000");
    gpmc_send('1',x"2772",x"3D03");
    gpmc_send('1',x"2773",x"0000");
    gpmc_send('1',x"2774",x"3C04");
    gpmc_send('1',x"2775",x"0000");
    gpmc_send('1',x"2776",x"3B05");
    gpmc_send('1',x"2777",x"0000");
    gpmc_send('1',x"2778",x"3A06");
    gpmc_send('1',x"2779",x"0000");
    gpmc_send('1',x"277A",x"3907");
    gpmc_send('1',x"277B",x"0000");
    gpmc_send('1',x"277C",x"3808");
    gpmc_send('1',x"277D",x"0000");
    gpmc_send('1',x"277E",x"3709");
    gpmc_send('1',x"277F",x"0000");
    gpmc_send('1',x"2780",x"360A");
    gpmc_send('1',x"2781",x"0000");
    gpmc_send('1',x"2782",x"350B");
    gpmc_send('1',x"2783",x"0000");
    gpmc_send('1',x"2784",x"340C");
    gpmc_send('1',x"2785",x"0000");
    gpmc_send('1',x"2786",x"330D");
    gpmc_send('1',x"2787",x"0000");
    gpmc_send('1',x"2788",x"320E");
    gpmc_send('1',x"2789",x"0000");
    gpmc_send('1',x"278A",x"310F");
    gpmc_send('1',x"278B",x"0000");
    gpmc_send('1',x"278C",x"3010");
    gpmc_send('1',x"278D",x"0000");
    gpmc_send('1',x"278E",x"2F11");
    gpmc_send('1',x"278F",x"0000");
    gpmc_send('1',x"2790",x"2E12");
    gpmc_send('1',x"2791",x"0000");
    gpmc_send('1',x"2792",x"2D13");
    gpmc_send('1',x"2793",x"0000");
    gpmc_send('1',x"2794",x"2C14");
    gpmc_send('1',x"2795",x"0000");
    gpmc_send('1',x"2796",x"2B15");
    gpmc_send('1',x"2797",x"0000");
    gpmc_send('1',x"2798",x"2A16");
    gpmc_send('1',x"2799",x"0000");
    gpmc_send('1',x"279A",x"2917");
    gpmc_send('1',x"279B",x"0000");
    gpmc_send('1',x"279C",x"2818");
    gpmc_send('1',x"279D",x"0000");
    gpmc_send('1',x"279E",x"2719");
    gpmc_send('1',x"279F",x"0000");
    gpmc_send('1',x"27A0",x"261A");
    gpmc_send('1',x"27A1",x"0000");
    gpmc_send('1',x"27A2",x"251B");
    gpmc_send('1',x"27A3",x"0000");
    gpmc_send('1',x"27A4",x"241C");
    gpmc_send('1',x"27A5",x"0000");
    gpmc_send('1',x"27A6",x"231D");
    gpmc_send('1',x"27A7",x"0000");
    gpmc_send('1',x"27A8",x"221E");
    gpmc_send('1',x"27A9",x"0000");
    gpmc_send('1',x"27AA",x"211F");
    gpmc_send('1',x"27AB",x"0000");
    gpmc_send('1',x"27AC",x"2020");
    gpmc_send('1',x"27AD",x"0000");
    gpmc_send('1',x"27AE",x"1F21");
    gpmc_send('1',x"27AF",x"0000");
    gpmc_send('1',x"27B0",x"1E22");
    gpmc_send('1',x"27B1",x"0000");
    gpmc_send('1',x"27B2",x"1D23");
    gpmc_send('1',x"27B3",x"0000");
    gpmc_send('1',x"27B4",x"1C24");
    gpmc_send('1',x"27B5",x"0000");
    gpmc_send('1',x"27B6",x"1B25");
    gpmc_send('1',x"27B7",x"0000");
    gpmc_send('1',x"27B8",x"1A26");
    gpmc_send('1',x"27B9",x"0000");
    gpmc_send('1',x"27BA",x"1927");
    gpmc_send('1',x"27BB",x"0000");
    gpmc_send('1',x"27BC",x"1828");
    gpmc_send('1',x"27BD",x"0000");
    gpmc_send('1',x"27BE",x"1729");
    gpmc_send('1',x"27BF",x"0000");
    gpmc_send('1',x"27C0",x"162A");
    gpmc_send('1',x"27C1",x"0000");
    gpmc_send('1',x"27C2",x"152B");
    gpmc_send('1',x"27C3",x"0000");
    gpmc_send('1',x"27C4",x"142C");
    gpmc_send('1',x"27C5",x"0000");
    gpmc_send('1',x"27C6",x"132D");
    gpmc_send('1',x"27C7",x"0000");
    gpmc_send('1',x"27C8",x"122E");
    gpmc_send('1',x"27C9",x"0000");
    gpmc_send('1',x"27CA",x"112F");
    gpmc_send('1',x"27CB",x"0000");
    gpmc_send('1',x"27CC",x"1030");
    gpmc_send('1',x"27CD",x"0000");
    gpmc_send('1',x"27CE",x"0F31");
    gpmc_send('1',x"27CF",x"0000");
    gpmc_send('1',x"27D0",x"0E32");
    gpmc_send('1',x"27D1",x"0000");
    gpmc_send('1',x"27D2",x"0D33");
    gpmc_send('1',x"27D3",x"0000");
    gpmc_send('1',x"27D4",x"0C34");
    gpmc_send('1',x"27D5",x"0000");
    gpmc_send('1',x"27D6",x"0B35");
    gpmc_send('1',x"27D7",x"0000");
    gpmc_send('1',x"27D8",x"0A36");
    gpmc_send('1',x"27D9",x"0000");
    gpmc_send('1',x"27DA",x"0937");
    gpmc_send('1',x"27DB",x"0000");
    gpmc_send('1',x"27DC",x"0838");
    gpmc_send('1',x"27DD",x"0000");
    gpmc_send('1',x"27DE",x"0739");
    gpmc_send('1',x"27DF",x"0000");
    gpmc_send('1',x"27E0",x"063A");
    gpmc_send('1',x"27E1",x"0000");
    gpmc_send('1',x"27E2",x"053B");
    gpmc_send('1',x"27E3",x"0000");
    gpmc_send('1',x"27E4",x"043C");
    gpmc_send('1',x"27E5",x"0000");
    gpmc_send('1',x"27E6",x"033D");
    gpmc_send('1',x"27E7",x"0000");
    gpmc_send('1',x"27E8",x"023E");
    gpmc_send('1',x"27E9",x"0000");
    gpmc_send('1',x"27EA",x"013F");
    gpmc_send('1',x"27EB",x"0000");
    gpmc_send('1',x"27EC",x"003F");
    gpmc_send('1',x"27ED",x"0000");
    gpmc_send('1',x"27EE",x"003E");
    gpmc_send('1',x"27EF",x"0001");
    gpmc_send('1',x"27F0",x"003D");
    gpmc_send('1',x"27F1",x"0002");
    gpmc_send('1',x"27F2",x"003C");
    gpmc_send('1',x"27F3",x"0003");
    gpmc_send('1',x"27F4",x"003B");
    gpmc_send('1',x"27F5",x"0004");
    gpmc_send('1',x"27F6",x"003A");
    gpmc_send('1',x"27F7",x"0005");
    gpmc_send('1',x"27F8",x"0039");
    gpmc_send('1',x"27F9",x"0006");
    gpmc_send('1',x"27FA",x"0038");
    gpmc_send('1',x"27FB",x"0007");
    gpmc_send('1',x"27FC",x"0037");
    gpmc_send('1',x"27FD",x"0008");
    gpmc_send('1',x"27FE",x"0036");
    gpmc_send('1',x"27FF",x"0009");
    gpmc_send('1',x"2800",x"0035");
    gpmc_send('1',x"2801",x"000A");
    gpmc_send('1',x"2802",x"0034");
    gpmc_send('1',x"2803",x"000B");
    gpmc_send('1',x"2804",x"0033");
    gpmc_send('1',x"2805",x"000C");
    gpmc_send('1',x"2806",x"0032");
    gpmc_send('1',x"2807",x"000D");
    gpmc_send('1',x"2808",x"0031");
    gpmc_send('1',x"2809",x"000E");
    gpmc_send('1',x"280A",x"0030");
    gpmc_send('1',x"280B",x"000F");
    gpmc_send('1',x"280C",x"002F");
    gpmc_send('1',x"280D",x"0010");
    gpmc_send('1',x"280E",x"002E");
    gpmc_send('1',x"280F",x"0011");
    gpmc_send('1',x"2810",x"002D");
    gpmc_send('1',x"2811",x"0012");
    gpmc_send('1',x"2812",x"002C");
    gpmc_send('1',x"2813",x"0013");
    gpmc_send('1',x"2814",x"002B");
    gpmc_send('1',x"2815",x"0014");
    gpmc_send('1',x"2816",x"002A");
    gpmc_send('1',x"2817",x"0015");
    gpmc_send('1',x"2818",x"0029");
    gpmc_send('1',x"2819",x"0016");
    gpmc_send('1',x"281A",x"0028");
    gpmc_send('1',x"281B",x"0017");
    gpmc_send('1',x"281C",x"0027");
    gpmc_send('1',x"281D",x"0018");
    gpmc_send('1',x"281E",x"0026");
    gpmc_send('1',x"281F",x"0019");
    gpmc_send('1',x"2820",x"0025");
    gpmc_send('1',x"2821",x"001A");
    gpmc_send('1',x"2822",x"0024");
    gpmc_send('1',x"2823",x"001B");
    gpmc_send('1',x"2824",x"0023");
    gpmc_send('1',x"2825",x"001C");
    gpmc_send('1',x"2826",x"0022");
    gpmc_send('1',x"2827",x"001D");
    gpmc_send('1',x"2828",x"0021");
    gpmc_send('1',x"2829",x"001E");
    gpmc_send('1',x"282A",x"0020");
    gpmc_send('1',x"282B",x"001F");
    gpmc_send('1',x"282C",x"001F");
    gpmc_send('1',x"282D",x"0020");
    gpmc_send('1',x"282E",x"001E");
    gpmc_send('1',x"282F",x"0021");
    gpmc_send('1',x"2830",x"001D");
    gpmc_send('1',x"2831",x"0022");
    gpmc_send('1',x"2832",x"001C");
    gpmc_send('1',x"2833",x"0023");
    gpmc_send('1',x"2834",x"001B");
    gpmc_send('1',x"2835",x"0024");
    gpmc_send('1',x"2836",x"001A");
    gpmc_send('1',x"2837",x"0025");
    gpmc_send('1',x"2838",x"0019");
    gpmc_send('1',x"2839",x"0026");
    gpmc_send('1',x"283A",x"0018");
    gpmc_send('1',x"283B",x"0027");
    gpmc_send('1',x"283C",x"0017");
    gpmc_send('1',x"283D",x"0028");
    gpmc_send('1',x"283E",x"0016");
    gpmc_send('1',x"283F",x"0029");
    gpmc_send('1',x"2840",x"0015");
    gpmc_send('1',x"2841",x"002A");
    gpmc_send('1',x"2842",x"0014");
    gpmc_send('1',x"2843",x"002B");
    gpmc_send('1',x"2844",x"0013");
    gpmc_send('1',x"2845",x"002C");
    gpmc_send('1',x"2846",x"0012");
    gpmc_send('1',x"2847",x"002D");
    gpmc_send('1',x"2848",x"0011");
    gpmc_send('1',x"2849",x"002E");
    gpmc_send('1',x"284A",x"0010");
    gpmc_send('1',x"284B",x"002F");
    gpmc_send('1',x"284C",x"000F");
    gpmc_send('1',x"284D",x"0030");
    gpmc_send('1',x"284E",x"000E");
    gpmc_send('1',x"284F",x"0031");
    gpmc_send('1',x"2850",x"000D");
    gpmc_send('1',x"2851",x"0032");
    gpmc_send('1',x"2852",x"000C");
    gpmc_send('1',x"2853",x"0033");
    gpmc_send('1',x"2854",x"000B");
    gpmc_send('1',x"2855",x"0034");
    gpmc_send('1',x"2856",x"000A");
    gpmc_send('1',x"2857",x"0035");
    gpmc_send('1',x"2858",x"0009");
    gpmc_send('1',x"2859",x"0036");
    gpmc_send('1',x"285A",x"0008");
    gpmc_send('1',x"285B",x"0037");
    gpmc_send('1',x"285C",x"0007");
    gpmc_send('1',x"285D",x"0038");
    gpmc_send('1',x"285E",x"0006");
    gpmc_send('1',x"285F",x"0039");
    gpmc_send('1',x"2860",x"0005");
    gpmc_send('1',x"2861",x"003A");
    gpmc_send('1',x"2862",x"0004");
    gpmc_send('1',x"2863",x"003B");
    gpmc_send('1',x"2864",x"0003");
    gpmc_send('1',x"2865",x"003C");
    gpmc_send('1',x"2866",x"0002");
    gpmc_send('1',x"2867",x"003D");
    gpmc_send('1',x"2868",x"0001");
    gpmc_send('1',x"2869",x"003E");
    gpmc_send('1',x"286A",x"0000");
    gpmc_send('1',x"286B",x"003F");
    gpmc_send('1',x"286C",x"0100");
    gpmc_send('1',x"286D",x"003E");
    gpmc_send('1',x"286E",x"0200");
    gpmc_send('1',x"286F",x"003D");
    gpmc_send('1',x"2870",x"0300");
    gpmc_send('1',x"2871",x"003C");
    gpmc_send('1',x"2872",x"0400");
    gpmc_send('1',x"2873",x"003B");
    gpmc_send('1',x"2874",x"0500");
    gpmc_send('1',x"2875",x"003A");
    gpmc_send('1',x"2876",x"0600");
    gpmc_send('1',x"2877",x"0039");
    gpmc_send('1',x"2878",x"0700");
    gpmc_send('1',x"2879",x"0038");
    gpmc_send('1',x"287A",x"0800");
    gpmc_send('1',x"287B",x"0037");
    gpmc_send('1',x"287C",x"0900");
    gpmc_send('1',x"287D",x"0036");
    gpmc_send('1',x"287E",x"0A00");
    gpmc_send('1',x"287F",x"0035");
    gpmc_send('1',x"2880",x"0B00");
    gpmc_send('1',x"2881",x"0034");
    gpmc_send('1',x"2882",x"0C00");
    gpmc_send('1',x"2883",x"0033");
    gpmc_send('1',x"2884",x"0D00");
    gpmc_send('1',x"2885",x"0032");
    gpmc_send('1',x"2886",x"0E00");
    gpmc_send('1',x"2887",x"0031");
    gpmc_send('1',x"2888",x"0F00");
    gpmc_send('1',x"2889",x"0030");
    gpmc_send('1',x"288A",x"1000");
    gpmc_send('1',x"288B",x"002F");
    gpmc_send('1',x"288C",x"1100");
    gpmc_send('1',x"288D",x"002E");
    gpmc_send('1',x"288E",x"1200");
    gpmc_send('1',x"288F",x"002D");
    gpmc_send('1',x"2890",x"1300");
    gpmc_send('1',x"2891",x"002C");
    gpmc_send('1',x"2892",x"1400");
    gpmc_send('1',x"2893",x"002B");
    gpmc_send('1',x"2894",x"1500");
    gpmc_send('1',x"2895",x"002A");
    gpmc_send('1',x"2896",x"1600");
    gpmc_send('1',x"2897",x"0029");
    gpmc_send('1',x"2898",x"1700");
    gpmc_send('1',x"2899",x"0028");
    gpmc_send('1',x"289A",x"1800");
    gpmc_send('1',x"289B",x"0027");
    gpmc_send('1',x"289C",x"1900");
    gpmc_send('1',x"289D",x"0026");
    gpmc_send('1',x"289E",x"1A00");
    gpmc_send('1',x"289F",x"0025");
    gpmc_send('1',x"28A0",x"1B00");
    gpmc_send('1',x"28A1",x"0024");
    gpmc_send('1',x"28A2",x"1C00");
    gpmc_send('1',x"28A3",x"0023");
    gpmc_send('1',x"28A4",x"1D00");
    gpmc_send('1',x"28A5",x"0022");
    gpmc_send('1',x"28A6",x"1E00");
    gpmc_send('1',x"28A7",x"0021");
    gpmc_send('1',x"28A8",x"1F00");
    gpmc_send('1',x"28A9",x"0020");
    gpmc_send('1',x"28AA",x"2000");
    gpmc_send('1',x"28AB",x"001F");
    gpmc_send('1',x"28AC",x"2100");
    gpmc_send('1',x"28AD",x"001E");
    gpmc_send('1',x"28AE",x"2200");
    gpmc_send('1',x"28AF",x"001D");
    gpmc_send('1',x"28B0",x"2300");
    gpmc_send('1',x"28B1",x"001C");
    gpmc_send('1',x"28B2",x"2400");
    gpmc_send('1',x"28B3",x"001B");
    gpmc_send('1',x"28B4",x"2500");
    gpmc_send('1',x"28B5",x"001A");
    gpmc_send('1',x"28B6",x"2600");
    gpmc_send('1',x"28B7",x"0019");
    gpmc_send('1',x"28B8",x"2700");
    gpmc_send('1',x"28B9",x"0018");
    gpmc_send('1',x"28BA",x"2800");
    gpmc_send('1',x"28BB",x"0017");
    gpmc_send('1',x"28BC",x"2900");
    gpmc_send('1',x"28BD",x"0016");
    gpmc_send('1',x"28BE",x"2A00");
    gpmc_send('1',x"28BF",x"0015");
    gpmc_send('1',x"28C0",x"2B00");
    gpmc_send('1',x"28C1",x"0014");
    gpmc_send('1',x"28C2",x"2C00");
    gpmc_send('1',x"28C3",x"0013");
    gpmc_send('1',x"28C4",x"2D00");
    gpmc_send('1',x"28C5",x"0012");
    gpmc_send('1',x"28C6",x"2E00");
    gpmc_send('1',x"28C7",x"0011");
    gpmc_send('1',x"28C8",x"2F00");
    gpmc_send('1',x"28C9",x"0010");
    gpmc_send('1',x"28CA",x"3000");
    gpmc_send('1',x"28CB",x"000F");
    gpmc_send('1',x"28CC",x"3100");
    gpmc_send('1',x"28CD",x"000E");
    gpmc_send('1',x"28CE",x"3200");
    gpmc_send('1',x"28CF",x"000D");
    gpmc_send('1',x"28D0",x"3300");
    gpmc_send('1',x"28D1",x"000C");
    gpmc_send('1',x"28D2",x"3400");
    gpmc_send('1',x"28D3",x"000B");
    gpmc_send('1',x"28D4",x"3500");
    gpmc_send('1',x"28D5",x"000A");
    gpmc_send('1',x"28D6",x"3600");
    gpmc_send('1',x"28D7",x"0009");
    gpmc_send('1',x"28D8",x"3700");
    gpmc_send('1',x"28D9",x"0008");
    gpmc_send('1',x"28DA",x"3800");
    gpmc_send('1',x"28DB",x"0007");
    gpmc_send('1',x"28DC",x"3900");
    gpmc_send('1',x"28DD",x"0006");
    gpmc_send('1',x"28DE",x"3A00");
    gpmc_send('1',x"28DF",x"0005");
    gpmc_send('1',x"28E0",x"3B00");
    gpmc_send('1',x"28E1",x"0004");
    gpmc_send('1',x"28E2",x"3C00");
    gpmc_send('1',x"28E3",x"0003");
    gpmc_send('1',x"28E4",x"3D00");
    gpmc_send('1',x"28E5",x"0002");
    gpmc_send('1',x"28E6",x"3E00");
    gpmc_send('1',x"28E7",x"0001");
    gpmc_send('1',x"28E8",x"3F00");
    gpmc_send('1',x"28E9",x"0000");
    gpmc_send('1',x"28EA",x"3F01");
    gpmc_send('1',x"28EB",x"0000");
    gpmc_send('1',x"28EC",x"3E02");
    gpmc_send('1',x"28ED",x"0000");
    gpmc_send('1',x"28EE",x"3D03");
    gpmc_send('1',x"28EF",x"0000");
    gpmc_send('1',x"28F0",x"3C04");
    gpmc_send('1',x"28F1",x"0000");
    gpmc_send('1',x"28F2",x"3B05");
    gpmc_send('1',x"28F3",x"0000");
    gpmc_send('1',x"28F4",x"3A06");
    gpmc_send('1',x"28F5",x"0000");
    gpmc_send('1',x"28F6",x"3907");
    gpmc_send('1',x"28F7",x"0000");
    gpmc_send('1',x"28F8",x"3808");
    gpmc_send('1',x"28F9",x"0000");
    gpmc_send('1',x"28FA",x"3709");
    gpmc_send('1',x"28FB",x"0000");
    gpmc_send('1',x"28FC",x"360A");
    gpmc_send('1',x"28FD",x"0000");
    gpmc_send('1',x"28FE",x"350B");
    gpmc_send('1',x"28FF",x"0000");
    gpmc_send('1',x"2900",x"340C");
    gpmc_send('1',x"2901",x"0000");
    gpmc_send('1',x"2902",x"330D");
    gpmc_send('1',x"2903",x"0000");
    gpmc_send('1',x"2904",x"320E");
    gpmc_send('1',x"2905",x"0000");
    gpmc_send('1',x"2906",x"310F");
    gpmc_send('1',x"2907",x"0000");
    gpmc_send('1',x"2908",x"3010");
    gpmc_send('1',x"2909",x"0000");
    gpmc_send('1',x"290A",x"2F11");
    gpmc_send('1',x"290B",x"0000");
    gpmc_send('1',x"290C",x"2E12");
    gpmc_send('1',x"290D",x"0000");
    gpmc_send('1',x"290E",x"2D13");
    gpmc_send('1',x"290F",x"0000");
    gpmc_send('1',x"2910",x"2C14");
    gpmc_send('1',x"2911",x"0000");
    gpmc_send('1',x"2912",x"2B15");
    gpmc_send('1',x"2913",x"0000");
    gpmc_send('1',x"2914",x"2A16");
    gpmc_send('1',x"2915",x"0000");
    gpmc_send('1',x"2916",x"2917");
    gpmc_send('1',x"2917",x"0000");
    gpmc_send('1',x"2918",x"2818");
    gpmc_send('1',x"2919",x"0000");
    gpmc_send('1',x"291A",x"2719");
    gpmc_send('1',x"291B",x"0000");
    gpmc_send('1',x"291C",x"261A");
    gpmc_send('1',x"291D",x"0000");
    gpmc_send('1',x"291E",x"251B");
    gpmc_send('1',x"291F",x"0000");
    gpmc_send('1',x"2920",x"241C");
    gpmc_send('1',x"2921",x"0000");
    gpmc_send('1',x"2922",x"231D");
    gpmc_send('1',x"2923",x"0000");
    gpmc_send('1',x"2924",x"221E");
    gpmc_send('1',x"2925",x"0000");
    gpmc_send('1',x"2926",x"211F");
    gpmc_send('1',x"2927",x"0000");
    gpmc_send('1',x"2928",x"2020");
    gpmc_send('1',x"2929",x"0000");
    gpmc_send('1',x"292A",x"1F21");
    gpmc_send('1',x"292B",x"0000");
    gpmc_send('1',x"292C",x"1E22");
    gpmc_send('1',x"292D",x"0000");
    gpmc_send('1',x"292E",x"1D23");
    gpmc_send('1',x"292F",x"0000");
    gpmc_send('1',x"2930",x"1C24");
    gpmc_send('1',x"2931",x"0000");
    gpmc_send('1',x"2932",x"1B25");
    gpmc_send('1',x"2933",x"0000");
    gpmc_send('1',x"2934",x"1A26");
    gpmc_send('1',x"2935",x"0000");
    gpmc_send('1',x"2936",x"1927");
    gpmc_send('1',x"2937",x"0000");
    gpmc_send('1',x"2938",x"1828");
    gpmc_send('1',x"2939",x"0000");
    gpmc_send('1',x"293A",x"1729");
    gpmc_send('1',x"293B",x"0000");
    gpmc_send('1',x"293C",x"162A");
    gpmc_send('1',x"293D",x"0000");
    gpmc_send('1',x"293E",x"152B");
    gpmc_send('1',x"293F",x"0000");
    gpmc_send('1',x"2940",x"142C");
    gpmc_send('1',x"2941",x"0000");
    gpmc_send('1',x"2942",x"132D");
    gpmc_send('1',x"2943",x"0000");
    gpmc_send('1',x"2944",x"122E");
    gpmc_send('1',x"2945",x"0000");
    gpmc_send('1',x"2946",x"112F");
    gpmc_send('1',x"2947",x"0000");
    gpmc_send('1',x"2948",x"1030");
    gpmc_send('1',x"2949",x"0000");
    gpmc_send('1',x"294A",x"0F31");
    gpmc_send('1',x"294B",x"0000");
    gpmc_send('1',x"294C",x"0E32");
    gpmc_send('1',x"294D",x"0000");
    gpmc_send('1',x"294E",x"0D33");
    gpmc_send('1',x"294F",x"0000");
    gpmc_send('1',x"2950",x"0C34");
    gpmc_send('1',x"2951",x"0000");
    gpmc_send('1',x"2952",x"0B35");
    gpmc_send('1',x"2953",x"0000");
    gpmc_send('1',x"2954",x"0A36");
    gpmc_send('1',x"2955",x"0000");
    gpmc_send('1',x"2956",x"0937");
    gpmc_send('1',x"2957",x"0000");
    gpmc_send('1',x"2958",x"0838");
    gpmc_send('1',x"2959",x"0000");
    gpmc_send('1',x"295A",x"0739");
    gpmc_send('1',x"295B",x"0000");
    gpmc_send('1',x"295C",x"063A");
    gpmc_send('1',x"295D",x"0000");
    gpmc_send('1',x"295E",x"053B");
    gpmc_send('1',x"295F",x"0000");
    gpmc_send('1',x"2960",x"043C");
    gpmc_send('1',x"2961",x"0000");
    gpmc_send('1',x"2962",x"033D");
    gpmc_send('1',x"2963",x"0000");
    gpmc_send('1',x"2964",x"023E");
    gpmc_send('1',x"2965",x"0000");
    gpmc_send('1',x"2966",x"013F");
    gpmc_send('1',x"2967",x"0000");
    gpmc_send('1',x"2968",x"003F");
    gpmc_send('1',x"2969",x"0000");
    gpmc_send('1',x"296A",x"003E");
    gpmc_send('1',x"296B",x"0001");
    gpmc_send('1',x"296C",x"003D");
    gpmc_send('1',x"296D",x"0002");
    gpmc_send('1',x"296E",x"003C");
    gpmc_send('1',x"296F",x"0003");
    gpmc_send('1',x"2970",x"003B");
    gpmc_send('1',x"2971",x"0004");
    gpmc_send('1',x"2972",x"003A");
    gpmc_send('1',x"2973",x"0005");
    gpmc_send('1',x"2974",x"0039");
    gpmc_send('1',x"2975",x"0006");
    gpmc_send('1',x"2976",x"0038");
    gpmc_send('1',x"2977",x"0007");
    gpmc_send('1',x"2978",x"0037");
    gpmc_send('1',x"2979",x"0008");
    gpmc_send('1',x"297A",x"0036");
    gpmc_send('1',x"297B",x"0009");
    gpmc_send('1',x"297C",x"0035");
    gpmc_send('1',x"297D",x"000A");
    gpmc_send('1',x"297E",x"0034");
    gpmc_send('1',x"297F",x"000B");
    gpmc_send('1',x"2980",x"0033");
    gpmc_send('1',x"2981",x"000C");
    gpmc_send('1',x"2982",x"0032");
    gpmc_send('1',x"2983",x"000D");
    gpmc_send('1',x"2984",x"0031");
    gpmc_send('1',x"2985",x"000E");
    gpmc_send('1',x"2986",x"0030");
    gpmc_send('1',x"2987",x"000F");
    gpmc_send('1',x"2988",x"002F");
    gpmc_send('1',x"2989",x"0010");
    gpmc_send('1',x"298A",x"002E");
    gpmc_send('1',x"298B",x"0011");
    gpmc_send('1',x"298C",x"002D");
    gpmc_send('1',x"298D",x"0012");
    gpmc_send('1',x"298E",x"002C");
    gpmc_send('1',x"298F",x"0013");
    gpmc_send('1',x"2990",x"002B");
    gpmc_send('1',x"2991",x"0014");
    gpmc_send('1',x"2992",x"002A");
    gpmc_send('1',x"2993",x"0015");
    gpmc_send('1',x"2994",x"0029");
    gpmc_send('1',x"2995",x"0016");
    gpmc_send('1',x"2996",x"0028");
    gpmc_send('1',x"2997",x"0017");
    gpmc_send('1',x"2998",x"0027");
    gpmc_send('1',x"2999",x"0018");
    gpmc_send('1',x"299A",x"0026");
    gpmc_send('1',x"299B",x"0019");
    gpmc_send('1',x"299C",x"0025");
    gpmc_send('1',x"299D",x"001A");
    gpmc_send('1',x"299E",x"0024");
    gpmc_send('1',x"299F",x"001B");
    gpmc_send('1',x"29A0",x"0023");
    gpmc_send('1',x"29A1",x"001C");
    gpmc_send('1',x"29A2",x"0022");
    gpmc_send('1',x"29A3",x"001D");
    gpmc_send('1',x"29A4",x"0021");
    gpmc_send('1',x"29A5",x"001E");
    gpmc_send('1',x"29A6",x"0020");
    gpmc_send('1',x"29A7",x"001F");
    gpmc_send('1',x"29A8",x"001F");
    gpmc_send('1',x"29A9",x"0020");
    gpmc_send('1',x"29AA",x"001E");
    gpmc_send('1',x"29AB",x"0021");
    gpmc_send('1',x"29AC",x"001D");
    gpmc_send('1',x"29AD",x"0022");
    gpmc_send('1',x"29AE",x"001C");
    gpmc_send('1',x"29AF",x"0023");
    gpmc_send('1',x"29B0",x"001B");
    gpmc_send('1',x"29B1",x"0024");
    gpmc_send('1',x"29B2",x"001A");
    gpmc_send('1',x"29B3",x"0025");
    gpmc_send('1',x"29B4",x"0019");
    gpmc_send('1',x"29B5",x"0026");
    gpmc_send('1',x"29B6",x"0018");
    gpmc_send('1',x"29B7",x"0027");
    gpmc_send('1',x"29B8",x"0017");
    gpmc_send('1',x"29B9",x"0028");
    gpmc_send('1',x"29BA",x"0016");
    gpmc_send('1',x"29BB",x"0029");
    gpmc_send('1',x"29BC",x"0015");
    gpmc_send('1',x"29BD",x"002A");
    gpmc_send('1',x"29BE",x"0014");
    gpmc_send('1',x"29BF",x"002B");
    gpmc_send('1',x"29C0",x"0013");
    gpmc_send('1',x"29C1",x"002C");
    gpmc_send('1',x"29C2",x"0012");
    gpmc_send('1',x"29C3",x"002D");
    gpmc_send('1',x"29C4",x"0011");
    gpmc_send('1',x"29C5",x"002E");
    gpmc_send('1',x"29C6",x"0010");
    gpmc_send('1',x"29C7",x"002F");
    gpmc_send('1',x"29C8",x"000F");
    gpmc_send('1',x"29C9",x"0030");
    gpmc_send('1',x"29CA",x"000E");
    gpmc_send('1',x"29CB",x"0031");
    gpmc_send('1',x"29CC",x"000D");
    gpmc_send('1',x"29CD",x"0032");
    gpmc_send('1',x"29CE",x"000C");
    gpmc_send('1',x"29CF",x"0033");
    gpmc_send('1',x"29D0",x"000B");
    gpmc_send('1',x"29D1",x"0034");
    gpmc_send('1',x"29D2",x"000A");
    gpmc_send('1',x"29D3",x"0035");
    gpmc_send('1',x"29D4",x"0009");
    gpmc_send('1',x"29D5",x"0036");
    gpmc_send('1',x"29D6",x"0008");
    gpmc_send('1',x"29D7",x"0037");
    gpmc_send('1',x"29D8",x"0007");
    gpmc_send('1',x"29D9",x"0038");
    gpmc_send('1',x"29DA",x"0006");
    gpmc_send('1',x"29DB",x"0039");
    gpmc_send('1',x"29DC",x"0005");
    gpmc_send('1',x"29DD",x"003A");
    gpmc_send('1',x"29DE",x"0004");
    gpmc_send('1',x"29DF",x"003B");
    gpmc_send('1',x"29E0",x"0003");
    gpmc_send('1',x"29E1",x"003C");
    gpmc_send('1',x"29E2",x"0002");
    gpmc_send('1',x"29E3",x"003D");
    gpmc_send('1',x"29E4",x"0001");
    gpmc_send('1',x"29E5",x"003E");
    gpmc_send('1',x"29E6",x"0000");
    gpmc_send('1',x"29E7",x"003F");
    gpmc_send('1',x"29E8",x"0100");
    gpmc_send('1',x"29E9",x"003E");
    gpmc_send('1',x"29EA",x"0200");
    gpmc_send('1',x"29EB",x"003D");
    gpmc_send('1',x"29EC",x"0300");
    gpmc_send('1',x"29ED",x"003C");
    gpmc_send('1',x"29EE",x"0400");
    gpmc_send('1',x"29EF",x"003B");
    gpmc_send('1',x"29F0",x"0500");
    gpmc_send('1',x"29F1",x"003A");
    gpmc_send('1',x"29F2",x"0600");
    gpmc_send('1',x"29F3",x"0039");
    gpmc_send('1',x"29F4",x"0700");
    gpmc_send('1',x"29F5",x"0038");
    gpmc_send('1',x"29F6",x"0800");
    gpmc_send('1',x"29F7",x"0037");
    gpmc_send('1',x"29F8",x"0900");
    gpmc_send('1',x"29F9",x"0036");
    gpmc_send('1',x"29FA",x"0A00");
    gpmc_send('1',x"29FB",x"0035");
    gpmc_send('1',x"29FC",x"0B00");
    gpmc_send('1',x"29FD",x"0034");
    gpmc_send('1',x"29FE",x"0C00");
    gpmc_send('1',x"29FF",x"0033");
    gpmc_send('1',x"2A00",x"0D00");
    gpmc_send('1',x"2A01",x"0032");
    gpmc_send('1',x"2A02",x"0E00");
    gpmc_send('1',x"2A03",x"0031");
    gpmc_send('1',x"2A04",x"0F00");
    gpmc_send('1',x"2A05",x"0030");
    gpmc_send('1',x"2A06",x"1000");
    gpmc_send('1',x"2A07",x"002F");
    gpmc_send('1',x"2A08",x"1100");
    gpmc_send('1',x"2A09",x"002E");
    gpmc_send('1',x"2A0A",x"1200");
    gpmc_send('1',x"2A0B",x"002D");
    gpmc_send('1',x"2A0C",x"1300");
    gpmc_send('1',x"2A0D",x"002C");
    gpmc_send('1',x"2A0E",x"1400");
    gpmc_send('1',x"2A0F",x"002B");
    gpmc_send('1',x"2A10",x"1500");
    gpmc_send('1',x"2A11",x"002A");
    gpmc_send('1',x"2A12",x"1600");
    gpmc_send('1',x"2A13",x"0029");
    gpmc_send('1',x"2A14",x"1700");
    gpmc_send('1',x"2A15",x"0028");
    gpmc_send('1',x"2A16",x"1800");
    gpmc_send('1',x"2A17",x"0027");
    gpmc_send('1',x"2A18",x"1900");
    gpmc_send('1',x"2A19",x"0026");
    gpmc_send('1',x"2A1A",x"1A00");
    gpmc_send('1',x"2A1B",x"0025");
    gpmc_send('1',x"2A1C",x"1B00");
    gpmc_send('1',x"2A1D",x"0024");
    gpmc_send('1',x"2A1E",x"1C00");
    gpmc_send('1',x"2A1F",x"0023");
    gpmc_send('1',x"2A20",x"1D00");
    gpmc_send('1',x"2A21",x"0022");
    gpmc_send('1',x"2A22",x"1E00");
    gpmc_send('1',x"2A23",x"0021");
    gpmc_send('1',x"2A24",x"1F00");
    gpmc_send('1',x"2A25",x"0020");
    gpmc_send('1',x"2A26",x"2000");
    gpmc_send('1',x"2A27",x"001F");
    gpmc_send('1',x"2A28",x"2100");
    gpmc_send('1',x"2A29",x"001E");
    gpmc_send('1',x"2A2A",x"2200");
    gpmc_send('1',x"2A2B",x"001D");
    gpmc_send('1',x"2A2C",x"2300");
    gpmc_send('1',x"2A2D",x"001C");
    gpmc_send('1',x"2A2E",x"2400");
    gpmc_send('1',x"2A2F",x"001B");
    gpmc_send('1',x"2A30",x"2500");
    gpmc_send('1',x"2A31",x"001A");
    gpmc_send('1',x"2A32",x"2600");
    gpmc_send('1',x"2A33",x"0019");
    gpmc_send('1',x"2A34",x"2700");
    gpmc_send('1',x"2A35",x"0018");
    gpmc_send('1',x"2A36",x"2800");
    gpmc_send('1',x"2A37",x"0017");
    gpmc_send('1',x"2A38",x"2900");
    gpmc_send('1',x"2A39",x"0016");
    gpmc_send('1',x"2A3A",x"2A00");
    gpmc_send('1',x"2A3B",x"0015");
    gpmc_send('1',x"2A3C",x"2B00");
    gpmc_send('1',x"2A3D",x"0014");
    gpmc_send('1',x"2A3E",x"2C00");
    gpmc_send('1',x"2A3F",x"0013");
    gpmc_send('1',x"2A40",x"2D00");
    gpmc_send('1',x"2A41",x"0012");
    gpmc_send('1',x"2A42",x"2E00");
    gpmc_send('1',x"2A43",x"0011");
    gpmc_send('1',x"2A44",x"2F00");
    gpmc_send('1',x"2A45",x"0010");
    gpmc_send('1',x"2A46",x"3000");
    gpmc_send('1',x"2A47",x"000F");
    gpmc_send('1',x"2A48",x"3100");
    gpmc_send('1',x"2A49",x"000E");
    gpmc_send('1',x"2A4A",x"3200");
    gpmc_send('1',x"2A4B",x"000D");
    gpmc_send('1',x"2A4C",x"3300");
    gpmc_send('1',x"2A4D",x"000C");
    gpmc_send('1',x"2A4E",x"3400");
    gpmc_send('1',x"2A4F",x"000B");
    gpmc_send('1',x"2A50",x"3500");
    gpmc_send('1',x"2A51",x"000A");
    gpmc_send('1',x"2A52",x"3600");
    gpmc_send('1',x"2A53",x"0009");
    gpmc_send('1',x"2A54",x"3700");
    gpmc_send('1',x"2A55",x"0008");
    gpmc_send('1',x"2A56",x"3800");
    gpmc_send('1',x"2A57",x"0007");
    gpmc_send('1',x"2A58",x"3900");
    gpmc_send('1',x"2A59",x"0006");
    gpmc_send('1',x"2A5A",x"3A00");
    gpmc_send('1',x"2A5B",x"0005");
    gpmc_send('1',x"2A5C",x"3B00");
    gpmc_send('1',x"2A5D",x"0004");
    gpmc_send('1',x"2A5E",x"3C00");
    gpmc_send('1',x"2A5F",x"0003");
    gpmc_send('1',x"2A60",x"3D00");
    gpmc_send('1',x"2A61",x"0002");
    gpmc_send('1',x"2A62",x"3E00");
    gpmc_send('1',x"2A63",x"0001");
    gpmc_send('1',x"2A64",x"3F00");
    gpmc_send('1',x"2A65",x"0000");
    gpmc_send('1',x"2A66",x"3F01");
    gpmc_send('1',x"2A67",x"0000");
    gpmc_send('1',x"2A68",x"3E02");
    gpmc_send('1',x"2A69",x"0000");
    gpmc_send('1',x"2A6A",x"3D03");
    gpmc_send('1',x"2A6B",x"0000");
    gpmc_send('1',x"2A6C",x"3C04");
    gpmc_send('1',x"2A6D",x"0000");
    gpmc_send('1',x"2A6E",x"3B05");
    gpmc_send('1',x"2A6F",x"0000");
    gpmc_send('1',x"2A70",x"3A06");
    gpmc_send('1',x"2A71",x"0000");
    gpmc_send('1',x"2A72",x"3907");
    gpmc_send('1',x"2A73",x"0000");
    gpmc_send('1',x"2A74",x"3808");
    gpmc_send('1',x"2A75",x"0000");
    gpmc_send('1',x"2A76",x"3709");
    gpmc_send('1',x"2A77",x"0000");
    gpmc_send('1',x"2A78",x"360A");
    gpmc_send('1',x"2A79",x"0000");
    gpmc_send('1',x"2A7A",x"350B");
    gpmc_send('1',x"2A7B",x"0000");
    gpmc_send('1',x"2A7C",x"340C");
    gpmc_send('1',x"2A7D",x"0000");
    gpmc_send('1',x"2A7E",x"330D");
    gpmc_send('1',x"2A7F",x"0000");
    gpmc_send('1',x"2A80",x"320E");
    gpmc_send('1',x"2A81",x"0000");
    gpmc_send('1',x"2A82",x"310F");
    gpmc_send('1',x"2A83",x"0000");
    gpmc_send('1',x"2A84",x"3010");
    gpmc_send('1',x"2A85",x"0000");
    gpmc_send('1',x"2A86",x"2F11");
    gpmc_send('1',x"2A87",x"0000");
    gpmc_send('1',x"2A88",x"2E12");
    gpmc_send('1',x"2A89",x"0000");
    gpmc_send('1',x"2A8A",x"2D13");
    gpmc_send('1',x"2A8B",x"0000");
    gpmc_send('1',x"2A8C",x"2C14");
    gpmc_send('1',x"2A8D",x"0000");
    gpmc_send('1',x"2A8E",x"2B15");
    gpmc_send('1',x"2A8F",x"0000");
    gpmc_send('1',x"2A90",x"2A16");
    gpmc_send('1',x"2A91",x"0000");
    gpmc_send('1',x"2A92",x"2917");
    gpmc_send('1',x"2A93",x"0000");
    gpmc_send('1',x"2A94",x"2818");
    gpmc_send('1',x"2A95",x"0000");
    gpmc_send('1',x"2A96",x"2719");
    gpmc_send('1',x"2A97",x"0000");
    gpmc_send('1',x"2A98",x"261A");
    gpmc_send('1',x"2A99",x"0000");
    gpmc_send('1',x"2A9A",x"251B");
    gpmc_send('1',x"2A9B",x"0000");
    gpmc_send('1',x"2A9C",x"241C");
    gpmc_send('1',x"2A9D",x"0000");
    gpmc_send('1',x"2A9E",x"231D");
    gpmc_send('1',x"2A9F",x"0000");
    gpmc_send('1',x"2AA0",x"221E");
    gpmc_send('1',x"2AA1",x"0000");
    gpmc_send('1',x"2AA2",x"211F");
    gpmc_send('1',x"2AA3",x"0000");
    gpmc_send('1',x"2AA4",x"2020");
    gpmc_send('1',x"2AA5",x"0000");
    gpmc_send('1',x"2AA6",x"1F21");
    gpmc_send('1',x"2AA7",x"0000");
    gpmc_send('1',x"2AA8",x"1E22");
    gpmc_send('1',x"2AA9",x"0000");
    gpmc_send('1',x"2AAA",x"1D23");
    gpmc_send('1',x"2AAB",x"0000");
    gpmc_send('1',x"2AAC",x"1C24");
    gpmc_send('1',x"2AAD",x"0000");
    gpmc_send('1',x"2AAE",x"1B25");
    gpmc_send('1',x"2AAF",x"0000");
    gpmc_send('1',x"2AB0",x"1A26");
    gpmc_send('1',x"2AB1",x"0000");
    gpmc_send('1',x"2AB2",x"1927");
    gpmc_send('1',x"2AB3",x"0000");
    gpmc_send('1',x"2AB4",x"1828");
    gpmc_send('1',x"2AB5",x"0000");
    gpmc_send('1',x"2AB6",x"1729");
    gpmc_send('1',x"2AB7",x"0000");
    gpmc_send('1',x"2AB8",x"162A");
    gpmc_send('1',x"2AB9",x"0000");
    gpmc_send('1',x"2ABA",x"152B");
    gpmc_send('1',x"2ABB",x"0000");
    gpmc_send('1',x"2ABC",x"142C");
    gpmc_send('1',x"2ABD",x"0000");
    gpmc_send('1',x"2ABE",x"132D");
    gpmc_send('1',x"2ABF",x"0000");
    gpmc_send('1',x"2AC0",x"122E");
    gpmc_send('1',x"2AC1",x"0000");
    gpmc_send('1',x"2AC2",x"112F");
    gpmc_send('1',x"2AC3",x"0000");
    gpmc_send('1',x"2AC4",x"1030");
    gpmc_send('1',x"2AC5",x"0000");
    gpmc_send('1',x"2AC6",x"0F31");
    gpmc_send('1',x"2AC7",x"0000");
    gpmc_send('1',x"2AC8",x"0E32");
    gpmc_send('1',x"2AC9",x"0000");
    gpmc_send('1',x"2ACA",x"0D33");
    gpmc_send('1',x"2ACB",x"0000");
    gpmc_send('1',x"2ACC",x"0C34");
    gpmc_send('1',x"2ACD",x"0000");
    gpmc_send('1',x"2ACE",x"0B35");
    gpmc_send('1',x"2ACF",x"0000");
    gpmc_send('1',x"2AD0",x"0A36");
    gpmc_send('1',x"2AD1",x"0000");
    gpmc_send('1',x"2AD2",x"0937");
    gpmc_send('1',x"2AD3",x"0000");
    gpmc_send('1',x"2AD4",x"0838");
    gpmc_send('1',x"2AD5",x"0000");
    gpmc_send('1',x"2AD6",x"0739");
    gpmc_send('1',x"2AD7",x"0000");
    gpmc_send('1',x"2AD8",x"063A");
    gpmc_send('1',x"2AD9",x"0000");
    gpmc_send('1',x"2ADA",x"053B");
    gpmc_send('1',x"2ADB",x"0000");
    gpmc_send('1',x"2ADC",x"043C");
    gpmc_send('1',x"2ADD",x"0000");
    gpmc_send('1',x"2ADE",x"033D");
    gpmc_send('1',x"2ADF",x"0000");
    gpmc_send('1',x"2AE0",x"023E");
    gpmc_send('1',x"2AE1",x"0000");
    gpmc_send('1',x"2AE2",x"013F");
    gpmc_send('1',x"2AE3",x"0000");
    gpmc_send('1',x"2AE4",x"003F");
    gpmc_send('1',x"2AE5",x"0000");
    gpmc_send('1',x"2AE6",x"003E");
    gpmc_send('1',x"2AE7",x"0001");
    gpmc_send('1',x"2AE8",x"003D");
    gpmc_send('1',x"2AE9",x"0002");
    gpmc_send('1',x"2AEA",x"003C");
    gpmc_send('1',x"2AEB",x"0003");
    gpmc_send('1',x"2AEC",x"003B");
    gpmc_send('1',x"2AED",x"0004");
    gpmc_send('1',x"2AEE",x"003A");
    gpmc_send('1',x"2AEF",x"0005");
    gpmc_send('1',x"2AF0",x"0039");
    gpmc_send('1',x"2AF1",x"0006");
    gpmc_send('1',x"2AF2",x"0038");
    gpmc_send('1',x"2AF3",x"0007");
    gpmc_send('1',x"2AF4",x"0037");
    gpmc_send('1',x"2AF5",x"0008");
    gpmc_send('1',x"2AF6",x"0036");
    gpmc_send('1',x"2AF7",x"0009");
    gpmc_send('1',x"2AF8",x"0035");
    gpmc_send('1',x"2AF9",x"000A");
    gpmc_send('1',x"2AFA",x"0034");
    gpmc_send('1',x"2AFB",x"000B");
    gpmc_send('1',x"2AFC",x"0033");
    gpmc_send('1',x"2AFD",x"000C");
    gpmc_send('1',x"2AFE",x"0032");
    gpmc_send('1',x"2AFF",x"000D");
    gpmc_send('1',x"2B00",x"0031");
    gpmc_send('1',x"2B01",x"000E");
    gpmc_send('1',x"2B02",x"0030");
    gpmc_send('1',x"2B03",x"000F");
    gpmc_send('1',x"2B04",x"002F");
    gpmc_send('1',x"2B05",x"0010");
    gpmc_send('1',x"2B06",x"002E");
    gpmc_send('1',x"2B07",x"0011");
    gpmc_send('1',x"2B08",x"002D");
    gpmc_send('1',x"2B09",x"0012");
    gpmc_send('1',x"2B0A",x"002C");
    gpmc_send('1',x"2B0B",x"0013");
    gpmc_send('1',x"2B0C",x"002B");
    gpmc_send('1',x"2B0D",x"0014");
    gpmc_send('1',x"2B0E",x"002A");
    gpmc_send('1',x"2B0F",x"0015");
    gpmc_send('1',x"2B10",x"0029");
    gpmc_send('1',x"2B11",x"0016");
    gpmc_send('1',x"2B12",x"0028");
    gpmc_send('1',x"2B13",x"0017");
    gpmc_send('1',x"2B14",x"0027");
    gpmc_send('1',x"2B15",x"0018");
    gpmc_send('1',x"2B16",x"0026");
    gpmc_send('1',x"2B17",x"0019");
    gpmc_send('1',x"2B18",x"0025");
    gpmc_send('1',x"2B19",x"001A");
    gpmc_send('1',x"2B1A",x"0024");
    gpmc_send('1',x"2B1B",x"001B");
    gpmc_send('1',x"2B1C",x"0023");
    gpmc_send('1',x"2B1D",x"001C");
    gpmc_send('1',x"2B1E",x"0022");
    gpmc_send('1',x"2B1F",x"001D");
    gpmc_send('1',x"2B20",x"0021");
    gpmc_send('1',x"2B21",x"001E");
    gpmc_send('1',x"2B22",x"0020");
    gpmc_send('1',x"2B23",x"001F");
    gpmc_send('1',x"2B24",x"001F");
    gpmc_send('1',x"2B25",x"0020");
    gpmc_send('1',x"2B26",x"001E");
    gpmc_send('1',x"2B27",x"0021");
    gpmc_send('1',x"2B28",x"001D");
    gpmc_send('1',x"2B29",x"0022");
    gpmc_send('1',x"2B2A",x"001C");
    gpmc_send('1',x"2B2B",x"0023");
    gpmc_send('1',x"2B2C",x"001B");
    gpmc_send('1',x"2B2D",x"0024");
    gpmc_send('1',x"2B2E",x"001A");
    gpmc_send('1',x"2B2F",x"0025");
    gpmc_send('1',x"2B30",x"0019");
    gpmc_send('1',x"2B31",x"0026");
    gpmc_send('1',x"2B32",x"0018");
    gpmc_send('1',x"2B33",x"0027");
    gpmc_send('1',x"2B34",x"0017");
    gpmc_send('1',x"2B35",x"0028");
    gpmc_send('1',x"2B36",x"0016");
    gpmc_send('1',x"2B37",x"0029");
    gpmc_send('1',x"2B38",x"0015");
    gpmc_send('1',x"2B39",x"002A");
    gpmc_send('1',x"2B3A",x"0014");
    gpmc_send('1',x"2B3B",x"002B");
    gpmc_send('1',x"2B3C",x"0013");
    gpmc_send('1',x"2B3D",x"002C");
    gpmc_send('1',x"2B3E",x"0012");
    gpmc_send('1',x"2B3F",x"002D");
    gpmc_send('1',x"2B40",x"0011");
    gpmc_send('1',x"2B41",x"002E");
    gpmc_send('1',x"2B42",x"0010");
    gpmc_send('1',x"2B43",x"002F");
    gpmc_send('1',x"2B44",x"000F");
    gpmc_send('1',x"2B45",x"0030");
    gpmc_send('1',x"2B46",x"000E");
    gpmc_send('1',x"2B47",x"0031");
    gpmc_send('1',x"2B48",x"000D");
    gpmc_send('1',x"2B49",x"0032");
    gpmc_send('1',x"2B4A",x"000C");
    gpmc_send('1',x"2B4B",x"0033");
    gpmc_send('1',x"2B4C",x"000B");
    gpmc_send('1',x"2B4D",x"0034");
    gpmc_send('1',x"2B4E",x"000A");
    gpmc_send('1',x"2B4F",x"0035");
    gpmc_send('1',x"2B50",x"0009");
    gpmc_send('1',x"2B51",x"0036");
    gpmc_send('1',x"2B52",x"0008");
    gpmc_send('1',x"2B53",x"0037");
    gpmc_send('1',x"2B54",x"0007");
    gpmc_send('1',x"2B55",x"0038");
    gpmc_send('1',x"2B56",x"0006");
    gpmc_send('1',x"2B57",x"0039");
    gpmc_send('1',x"2B58",x"0005");
    gpmc_send('1',x"2B59",x"003A");
    gpmc_send('1',x"2B5A",x"0004");
    gpmc_send('1',x"2B5B",x"003B");
    gpmc_send('1',x"2B5C",x"0003");
    gpmc_send('1',x"2B5D",x"003C");
    gpmc_send('1',x"2B5E",x"0002");
    gpmc_send('1',x"2B5F",x"003D");
    gpmc_send('1',x"2B60",x"0001");
    gpmc_send('1',x"2B61",x"003E");
    gpmc_send('1',x"2B62",x"0000");
    gpmc_send('1',x"2B63",x"003F");
    gpmc_send('1',x"2B64",x"0100");
    gpmc_send('1',x"2B65",x"003E");
    gpmc_send('1',x"2B66",x"0200");
    gpmc_send('1',x"2B67",x"003D");
    gpmc_send('1',x"2B68",x"0300");
    gpmc_send('1',x"2B69",x"003C");
    gpmc_send('1',x"2B6A",x"0400");
    gpmc_send('1',x"2B6B",x"003B");
    gpmc_send('1',x"2B6C",x"0500");
    gpmc_send('1',x"2B6D",x"003A");
    gpmc_send('1',x"2B6E",x"0600");
    gpmc_send('1',x"2B6F",x"0039");
    gpmc_send('1',x"2B70",x"0700");
    gpmc_send('1',x"2B71",x"0038");
    gpmc_send('1',x"2B72",x"0800");
    gpmc_send('1',x"2B73",x"0037");
    gpmc_send('1',x"2B74",x"0900");
    gpmc_send('1',x"2B75",x"0036");
    gpmc_send('1',x"2B76",x"0A00");
    gpmc_send('1',x"2B77",x"0035");
    gpmc_send('1',x"2B78",x"0B00");
    gpmc_send('1',x"2B79",x"0034");
    gpmc_send('1',x"2B7A",x"0C00");
    gpmc_send('1',x"2B7B",x"0033");
    gpmc_send('1',x"2B7C",x"0D00");
    gpmc_send('1',x"2B7D",x"0032");
    gpmc_send('1',x"2B7E",x"0E00");
    gpmc_send('1',x"2B7F",x"0031");
    gpmc_send('1',x"2B80",x"0F00");
    gpmc_send('1',x"2B81",x"0030");
    gpmc_send('1',x"2B82",x"1000");
    gpmc_send('1',x"2B83",x"002F");
    gpmc_send('1',x"2B84",x"1100");
    gpmc_send('1',x"2B85",x"002E");
    gpmc_send('1',x"2B86",x"1200");
    gpmc_send('1',x"2B87",x"002D");
    gpmc_send('1',x"2B88",x"1300");
    gpmc_send('1',x"2B89",x"002C");
    gpmc_send('1',x"2B8A",x"1400");
    gpmc_send('1',x"2B8B",x"002B");
    gpmc_send('1',x"2B8C",x"1500");
    gpmc_send('1',x"2B8D",x"002A");
    gpmc_send('1',x"2B8E",x"1600");
    gpmc_send('1',x"2B8F",x"0029");
    gpmc_send('1',x"2B90",x"1700");
    gpmc_send('1',x"2B91",x"0028");
    gpmc_send('1',x"2B92",x"1800");
    gpmc_send('1',x"2B93",x"0027");
    gpmc_send('1',x"2B94",x"1900");
    gpmc_send('1',x"2B95",x"0026");
    gpmc_send('1',x"2B96",x"1A00");
    gpmc_send('1',x"2B97",x"0025");
    gpmc_send('1',x"2B98",x"1B00");
    gpmc_send('1',x"2B99",x"0024");
    gpmc_send('1',x"2B9A",x"1C00");
    gpmc_send('1',x"2B9B",x"0023");
    gpmc_send('1',x"2B9C",x"1D00");
    gpmc_send('1',x"2B9D",x"0022");
    gpmc_send('1',x"2B9E",x"1E00");
    gpmc_send('1',x"2B9F",x"0021");
    gpmc_send('1',x"2BA0",x"1F00");
    gpmc_send('1',x"2BA1",x"0020");
    gpmc_send('1',x"2BA2",x"2000");
    gpmc_send('1',x"2BA3",x"001F");
    gpmc_send('1',x"2BA4",x"2100");
    gpmc_send('1',x"2BA5",x"001E");
    gpmc_send('1',x"2BA6",x"2200");
    gpmc_send('1',x"2BA7",x"001D");
    gpmc_send('1',x"2BA8",x"2300");
    gpmc_send('1',x"2BA9",x"001C");
    gpmc_send('1',x"2BAA",x"2400");
    gpmc_send('1',x"2BAB",x"001B");
    gpmc_send('1',x"2BAC",x"2500");
    gpmc_send('1',x"2BAD",x"001A");
    gpmc_send('1',x"2BAE",x"2600");
    gpmc_send('1',x"2BAF",x"0019");
    gpmc_send('1',x"2BB0",x"2700");
    gpmc_send('1',x"2BB1",x"0018");
    gpmc_send('1',x"2BB2",x"2800");
    gpmc_send('1',x"2BB3",x"0017");
    gpmc_send('1',x"2BB4",x"2900");
    gpmc_send('1',x"2BB5",x"0016");
    gpmc_send('1',x"2BB6",x"2A00");
    gpmc_send('1',x"2BB7",x"0015");
    gpmc_send('1',x"2BB8",x"2B00");
    gpmc_send('1',x"2BB9",x"0014");
    gpmc_send('1',x"2BBA",x"2C00");
    gpmc_send('1',x"2BBB",x"0013");
    gpmc_send('1',x"2BBC",x"2D00");
    gpmc_send('1',x"2BBD",x"0012");
    gpmc_send('1',x"2BBE",x"2E00");
    gpmc_send('1',x"2BBF",x"0011");
    gpmc_send('1',x"2BC0",x"2F00");
    gpmc_send('1',x"2BC1",x"0010");
    gpmc_send('1',x"2BC2",x"3000");
    gpmc_send('1',x"2BC3",x"000F");
    gpmc_send('1',x"2BC4",x"3100");
    gpmc_send('1',x"2BC5",x"000E");
    gpmc_send('1',x"2BC6",x"3200");
    gpmc_send('1',x"2BC7",x"000D");
    gpmc_send('1',x"2BC8",x"3300");
    gpmc_send('1',x"2BC9",x"000C");
    gpmc_send('1',x"2BCA",x"3400");
    gpmc_send('1',x"2BCB",x"000B");
    gpmc_send('1',x"2BCC",x"3500");
    gpmc_send('1',x"2BCD",x"000A");
    gpmc_send('1',x"2BCE",x"3600");
    gpmc_send('1',x"2BCF",x"0009");
    gpmc_send('1',x"2BD0",x"3700");
    gpmc_send('1',x"2BD1",x"0008");
    gpmc_send('1',x"2BD2",x"3800");
    gpmc_send('1',x"2BD3",x"0007");
    gpmc_send('1',x"2BD4",x"3900");
    gpmc_send('1',x"2BD5",x"0006");
    gpmc_send('1',x"2BD6",x"3A00");
    gpmc_send('1',x"2BD7",x"0005");
    gpmc_send('1',x"2BD8",x"3B00");
    gpmc_send('1',x"2BD9",x"0004");
    gpmc_send('1',x"2BDA",x"3C00");
    gpmc_send('1',x"2BDB",x"0003");
    gpmc_send('1',x"2BDC",x"3D00");
    gpmc_send('1',x"2BDD",x"0002");
    gpmc_send('1',x"2BDE",x"3E00");
    gpmc_send('1',x"2BDF",x"0001");
    gpmc_send('1',x"2BE0",x"3F00");
    gpmc_send('1',x"2BE1",x"0000");
    gpmc_send('1',x"2BE2",x"3F01");
    gpmc_send('1',x"2BE3",x"0000");
    gpmc_send('1',x"2BE4",x"3E02");
    gpmc_send('1',x"2BE5",x"0000");
    gpmc_send('1',x"2BE6",x"3D03");
    gpmc_send('1',x"2BE7",x"0000");
    gpmc_send('1',x"2BE8",x"3C04");
    gpmc_send('1',x"2BE9",x"0000");
    gpmc_send('1',x"2BEA",x"3B05");
    gpmc_send('1',x"2BEB",x"0000");
    gpmc_send('1',x"2BEC",x"3A06");
    gpmc_send('1',x"2BED",x"0000");
    gpmc_send('1',x"2BEE",x"3907");
    gpmc_send('1',x"2BEF",x"0000");
    gpmc_send('1',x"2BF0",x"3808");
    gpmc_send('1',x"2BF1",x"0000");
    gpmc_send('1',x"2BF2",x"3709");
    gpmc_send('1',x"2BF3",x"0000");
    gpmc_send('1',x"2BF4",x"360A");
    gpmc_send('1',x"2BF5",x"0000");
    gpmc_send('1',x"2BF6",x"350B");
    gpmc_send('1',x"2BF7",x"0000");
    gpmc_send('1',x"2BF8",x"340C");
    gpmc_send('1',x"2BF9",x"0000");
    gpmc_send('1',x"2BFA",x"330D");
    gpmc_send('1',x"2BFB",x"0000");
    gpmc_send('1',x"2BFC",x"320E");
    gpmc_send('1',x"2BFD",x"0000");
    gpmc_send('1',x"2BFE",x"310F");
    gpmc_send('1',x"2BFF",x"0000");
    gpmc_send('1',x"2C00",x"3010");
    gpmc_send('1',x"2C01",x"0000");
    gpmc_send('1',x"2C02",x"2F11");
    gpmc_send('1',x"2C03",x"0000");
    gpmc_send('1',x"2C04",x"2E12");
    gpmc_send('1',x"2C05",x"0000");
    gpmc_send('1',x"2C06",x"2D13");
    gpmc_send('1',x"2C07",x"0000");
    gpmc_send('1',x"2C08",x"2C14");
    gpmc_send('1',x"2C09",x"0000");
    gpmc_send('1',x"2C0A",x"2B15");
    gpmc_send('1',x"2C0B",x"0000");
    gpmc_send('1',x"2C0C",x"2A16");
    gpmc_send('1',x"2C0D",x"0000");
    gpmc_send('1',x"2C0E",x"2917");
    gpmc_send('1',x"2C0F",x"0000");
    gpmc_send('1',x"2C10",x"2818");
    gpmc_send('1',x"2C11",x"0000");
    gpmc_send('1',x"2C12",x"2719");
    gpmc_send('1',x"2C13",x"0000");
    gpmc_send('1',x"2C14",x"261A");
    gpmc_send('1',x"2C15",x"0000");
    gpmc_send('1',x"2C16",x"251B");
    gpmc_send('1',x"2C17",x"0000");
    gpmc_send('1',x"2C18",x"241C");
    gpmc_send('1',x"2C19",x"0000");
    gpmc_send('1',x"2C1A",x"231D");
    gpmc_send('1',x"2C1B",x"0000");
    gpmc_send('1',x"2C1C",x"221E");
    gpmc_send('1',x"2C1D",x"0000");
    gpmc_send('1',x"2C1E",x"211F");
    gpmc_send('1',x"2C1F",x"0000");
    gpmc_send('1',x"2C20",x"2020");
    gpmc_send('1',x"2C21",x"0000");
    gpmc_send('1',x"2C22",x"1F21");
    gpmc_send('1',x"2C23",x"0000");
    gpmc_send('1',x"2C24",x"1E22");
    gpmc_send('1',x"2C25",x"0000");
    gpmc_send('1',x"2C26",x"1D23");
    gpmc_send('1',x"2C27",x"0000");
    gpmc_send('1',x"2C28",x"1C24");
    gpmc_send('1',x"2C29",x"0000");
    gpmc_send('1',x"2C2A",x"1B25");
    gpmc_send('1',x"2C2B",x"0000");
    gpmc_send('1',x"2C2C",x"1A26");
    gpmc_send('1',x"2C2D",x"0000");
    gpmc_send('1',x"2C2E",x"1927");
    gpmc_send('1',x"2C2F",x"0000");
    gpmc_send('1',x"2C30",x"1828");
    gpmc_send('1',x"2C31",x"0000");
    gpmc_send('1',x"2C32",x"1729");
    gpmc_send('1',x"2C33",x"0000");
    gpmc_send('1',x"2C34",x"162A");
    gpmc_send('1',x"2C35",x"0000");
    gpmc_send('1',x"2C36",x"152B");
    gpmc_send('1',x"2C37",x"0000");
    gpmc_send('1',x"2C38",x"142C");
    gpmc_send('1',x"2C39",x"0000");
    gpmc_send('1',x"2C3A",x"132D");
    gpmc_send('1',x"2C3B",x"0000");
    gpmc_send('1',x"2C3C",x"122E");
    gpmc_send('1',x"2C3D",x"0000");
    gpmc_send('1',x"2C3E",x"112F");
    gpmc_send('1',x"2C3F",x"0000");
    gpmc_send('1',x"2C40",x"1030");
    gpmc_send('1',x"2C41",x"0000");
    gpmc_send('1',x"2C42",x"0F31");
    gpmc_send('1',x"2C43",x"0000");
    gpmc_send('1',x"2C44",x"0E32");
    gpmc_send('1',x"2C45",x"0000");
    gpmc_send('1',x"2C46",x"0D33");
    gpmc_send('1',x"2C47",x"0000");
    gpmc_send('1',x"2C48",x"0C34");
    gpmc_send('1',x"2C49",x"0000");
    gpmc_send('1',x"2C4A",x"0B35");
    gpmc_send('1',x"2C4B",x"0000");
    gpmc_send('1',x"2C4C",x"0A36");
    gpmc_send('1',x"2C4D",x"0000");
    gpmc_send('1',x"2C4E",x"0937");
    gpmc_send('1',x"2C4F",x"0000");
    gpmc_send('1',x"2C50",x"0838");
    gpmc_send('1',x"2C51",x"0000");
    gpmc_send('1',x"2C52",x"0739");
    gpmc_send('1',x"2C53",x"0000");
    gpmc_send('1',x"2C54",x"063A");
    gpmc_send('1',x"2C55",x"0000");
    gpmc_send('1',x"2C56",x"053B");
    gpmc_send('1',x"2C57",x"0000");
    gpmc_send('1',x"2C58",x"043C");
    gpmc_send('1',x"2C59",x"0000");
    gpmc_send('1',x"2C5A",x"033D");
    gpmc_send('1',x"2C5B",x"0000");
    gpmc_send('1',x"2C5C",x"023E");
    gpmc_send('1',x"2C5D",x"0000");
    gpmc_send('1',x"2C5E",x"013F");
    gpmc_send('1',x"2C5F",x"0000");
    gpmc_send('1',x"2C60",x"003F");
    gpmc_send('1',x"2C61",x"0000");
    gpmc_send('1',x"2C62",x"003E");
    gpmc_send('1',x"2C63",x"0001");
    gpmc_send('1',x"2C64",x"003D");
    gpmc_send('1',x"2C65",x"0002");
    gpmc_send('1',x"2C66",x"003C");
    gpmc_send('1',x"2C67",x"0003");
    gpmc_send('1',x"2C68",x"003B");
    gpmc_send('1',x"2C69",x"0004");
    gpmc_send('1',x"2C6A",x"003A");
    gpmc_send('1',x"2C6B",x"0005");
    gpmc_send('1',x"2C6C",x"0039");
    gpmc_send('1',x"2C6D",x"0006");
    gpmc_send('1',x"2C6E",x"0038");
    gpmc_send('1',x"2C6F",x"0007");
    gpmc_send('1',x"2C70",x"0037");
    gpmc_send('1',x"2C71",x"0008");
    gpmc_send('1',x"2C72",x"0036");
    gpmc_send('1',x"2C73",x"0009");
    gpmc_send('1',x"2C74",x"0035");
    gpmc_send('1',x"2C75",x"000A");
    gpmc_send('1',x"2C76",x"0034");
    gpmc_send('1',x"2C77",x"000B");
    gpmc_send('1',x"2C78",x"0033");
    gpmc_send('1',x"2C79",x"000C");
    gpmc_send('1',x"2C7A",x"0032");
    gpmc_send('1',x"2C7B",x"000D");
    gpmc_send('1',x"2C7C",x"0031");
    gpmc_send('1',x"2C7D",x"000E");
    gpmc_send('1',x"2C7E",x"0030");
    gpmc_send('1',x"2C7F",x"000F");
    gpmc_send('1',x"2C80",x"002F");
    gpmc_send('1',x"2C81",x"0010");
    gpmc_send('1',x"2C82",x"002E");
    gpmc_send('1',x"2C83",x"0011");
    gpmc_send('1',x"2C84",x"002D");
    gpmc_send('1',x"2C85",x"0012");
    gpmc_send('1',x"2C86",x"002C");
    gpmc_send('1',x"2C87",x"0013");
    gpmc_send('1',x"2C88",x"002B");
    gpmc_send('1',x"2C89",x"0014");
    gpmc_send('1',x"2C8A",x"002A");
    gpmc_send('1',x"2C8B",x"0015");
    gpmc_send('1',x"2C8C",x"0029");
    gpmc_send('1',x"2C8D",x"0016");
    gpmc_send('1',x"2C8E",x"0028");
    gpmc_send('1',x"2C8F",x"0017");
    gpmc_send('1',x"2C90",x"0027");
    gpmc_send('1',x"2C91",x"0018");
    gpmc_send('1',x"2C92",x"0026");
    gpmc_send('1',x"2C93",x"0019");
    gpmc_send('1',x"2C94",x"0025");
    gpmc_send('1',x"2C95",x"001A");
    gpmc_send('1',x"2C96",x"0024");
    gpmc_send('1',x"2C97",x"001B");
    gpmc_send('1',x"2C98",x"0023");
    gpmc_send('1',x"2C99",x"001C");
    gpmc_send('1',x"2C9A",x"0022");
    gpmc_send('1',x"2C9B",x"001D");
    gpmc_send('1',x"2C9C",x"0021");
    gpmc_send('1',x"2C9D",x"001E");
    gpmc_send('1',x"2C9E",x"0020");
    gpmc_send('1',x"2C9F",x"001F");
    gpmc_send('1',x"2CA0",x"001F");
    gpmc_send('1',x"2CA1",x"0020");
    gpmc_send('1',x"2CA2",x"001E");
    gpmc_send('1',x"2CA3",x"0021");
    gpmc_send('1',x"2CA4",x"001D");
    gpmc_send('1',x"2CA5",x"0022");
    gpmc_send('1',x"2CA6",x"001C");
    gpmc_send('1',x"2CA7",x"0023");
    gpmc_send('1',x"2CA8",x"001B");
    gpmc_send('1',x"2CA9",x"0024");
    gpmc_send('1',x"2CAA",x"001A");
    gpmc_send('1',x"2CAB",x"0025");
    gpmc_send('1',x"2CAC",x"0019");
    gpmc_send('1',x"2CAD",x"0026");
    gpmc_send('1',x"2CAE",x"0018");
    gpmc_send('1',x"2CAF",x"0027");
    gpmc_send('1',x"2CB0",x"0017");
    gpmc_send('1',x"2CB1",x"0028");
    gpmc_send('1',x"2CB2",x"0016");
    gpmc_send('1',x"2CB3",x"0029");
    gpmc_send('1',x"2CB4",x"0015");
    gpmc_send('1',x"2CB5",x"002A");
    gpmc_send('1',x"2CB6",x"0014");
    gpmc_send('1',x"2CB7",x"002B");
    gpmc_send('1',x"2CB8",x"0013");
    gpmc_send('1',x"2CB9",x"002C");
    gpmc_send('1',x"2CBA",x"0012");
    gpmc_send('1',x"2CBB",x"002D");
    gpmc_send('1',x"2CBC",x"0011");
    gpmc_send('1',x"2CBD",x"002E");
    gpmc_send('1',x"2CBE",x"0010");
    gpmc_send('1',x"2CBF",x"002F");
    gpmc_send('1',x"2CC0",x"000F");
    gpmc_send('1',x"2CC1",x"0030");
    gpmc_send('1',x"2CC2",x"000E");
    gpmc_send('1',x"2CC3",x"0031");
    gpmc_send('1',x"2CC4",x"000D");
    gpmc_send('1',x"2CC5",x"0032");
    gpmc_send('1',x"2CC6",x"000C");
    gpmc_send('1',x"2CC7",x"0033");
    gpmc_send('1',x"2CC8",x"000B");
    gpmc_send('1',x"2CC9",x"0034");
    gpmc_send('1',x"2CCA",x"000A");
    gpmc_send('1',x"2CCB",x"0035");
    gpmc_send('1',x"2CCC",x"0009");
    gpmc_send('1',x"2CCD",x"0036");
    gpmc_send('1',x"2CCE",x"0008");
    gpmc_send('1',x"2CCF",x"0037");
    gpmc_send('1',x"2CD0",x"0007");
    gpmc_send('1',x"2CD1",x"0038");
    gpmc_send('1',x"2CD2",x"0006");
    gpmc_send('1',x"2CD3",x"0039");
    gpmc_send('1',x"2CD4",x"0005");
    gpmc_send('1',x"2CD5",x"003A");
    gpmc_send('1',x"2CD6",x"0004");
    gpmc_send('1',x"2CD7",x"003B");
    gpmc_send('1',x"2CD8",x"0003");
    gpmc_send('1',x"2CD9",x"003C");
    gpmc_send('1',x"2CDA",x"0002");
    gpmc_send('1',x"2CDB",x"003D");
    gpmc_send('1',x"2CDC",x"0001");
    gpmc_send('1',x"2CDD",x"003E");
    gpmc_send('1',x"2CDE",x"0000");
    gpmc_send('1',x"2CDF",x"003F");
    gpmc_send('1',x"2CE0",x"0100");
    gpmc_send('1',x"2CE1",x"003E");
    gpmc_send('1',x"2CE2",x"0200");
    gpmc_send('1',x"2CE3",x"003D");
    gpmc_send('1',x"2CE4",x"0300");
    gpmc_send('1',x"2CE5",x"003C");
    gpmc_send('1',x"2CE6",x"0400");
    gpmc_send('1',x"2CE7",x"003B");
    gpmc_send('1',x"2CE8",x"0500");
    gpmc_send('1',x"2CE9",x"003A");
    gpmc_send('1',x"2CEA",x"0600");
    gpmc_send('1',x"2CEB",x"0039");
    gpmc_send('1',x"2CEC",x"0700");
    gpmc_send('1',x"2CED",x"0038");
    gpmc_send('1',x"2CEE",x"0800");
    gpmc_send('1',x"2CEF",x"0037");
    gpmc_send('1',x"2CF0",x"0900");
    gpmc_send('1',x"2CF1",x"0036");
    gpmc_send('1',x"2CF2",x"0A00");
    gpmc_send('1',x"2CF3",x"0035");
    gpmc_send('1',x"2CF4",x"0B00");
    gpmc_send('1',x"2CF5",x"0034");
    gpmc_send('1',x"2CF6",x"0C00");
    gpmc_send('1',x"2CF7",x"0033");
    gpmc_send('1',x"2CF8",x"0D00");
    gpmc_send('1',x"2CF9",x"0032");
    gpmc_send('1',x"2CFA",x"0E00");
    gpmc_send('1',x"2CFB",x"0031");
    gpmc_send('1',x"2CFC",x"0F00");
    gpmc_send('1',x"2CFD",x"0030");
    gpmc_send('1',x"2CFE",x"1000");
    gpmc_send('1',x"2CFF",x"002F");
    gpmc_send('1',x"2D00",x"1100");
    gpmc_send('1',x"2D01",x"002E");
    gpmc_send('1',x"2D02",x"1200");
    gpmc_send('1',x"2D03",x"002D");
    gpmc_send('1',x"2D04",x"1300");
    gpmc_send('1',x"2D05",x"002C");
    gpmc_send('1',x"2D06",x"1400");
    gpmc_send('1',x"2D07",x"002B");
    gpmc_send('1',x"2D08",x"1500");
    gpmc_send('1',x"2D09",x"002A");
    gpmc_send('1',x"2D0A",x"1600");
    gpmc_send('1',x"2D0B",x"0029");
    gpmc_send('1',x"2D0C",x"1700");
    gpmc_send('1',x"2D0D",x"0028");
    gpmc_send('1',x"2D0E",x"1800");
    gpmc_send('1',x"2D0F",x"0027");
    gpmc_send('1',x"2D10",x"1900");
    gpmc_send('1',x"2D11",x"0026");
    gpmc_send('1',x"2D12",x"1A00");
    gpmc_send('1',x"2D13",x"0025");
    gpmc_send('1',x"2D14",x"1B00");
    gpmc_send('1',x"2D15",x"0024");
    gpmc_send('1',x"2D16",x"1C00");
    gpmc_send('1',x"2D17",x"0023");
    gpmc_send('1',x"2D18",x"1D00");
    gpmc_send('1',x"2D19",x"0022");
    gpmc_send('1',x"2D1A",x"1E00");
    gpmc_send('1',x"2D1B",x"0021");
    gpmc_send('1',x"2D1C",x"1F00");
    gpmc_send('1',x"2D1D",x"0020");
    gpmc_send('1',x"2D1E",x"2000");
    gpmc_send('1',x"2D1F",x"001F");
    gpmc_send('1',x"2D20",x"2100");
    gpmc_send('1',x"2D21",x"001E");
    gpmc_send('1',x"2D22",x"2200");
    gpmc_send('1',x"2D23",x"001D");
    gpmc_send('1',x"2D24",x"2300");
    gpmc_send('1',x"2D25",x"001C");
    gpmc_send('1',x"2D26",x"2400");
    gpmc_send('1',x"2D27",x"001B");
    gpmc_send('1',x"2D28",x"2500");
    gpmc_send('1',x"2D29",x"001A");
    gpmc_send('1',x"2D2A",x"2600");
    gpmc_send('1',x"2D2B",x"0019");
    gpmc_send('1',x"2D2C",x"2700");
    gpmc_send('1',x"2D2D",x"0018");
    gpmc_send('1',x"2D2E",x"2800");
    gpmc_send('1',x"2D2F",x"0017");
    gpmc_send('1',x"2D30",x"2900");
    gpmc_send('1',x"2D31",x"0016");
    gpmc_send('1',x"2D32",x"2A00");
    gpmc_send('1',x"2D33",x"0015");
    gpmc_send('1',x"2D34",x"2B00");
    gpmc_send('1',x"2D35",x"0014");
    gpmc_send('1',x"2D36",x"2C00");
    gpmc_send('1',x"2D37",x"0013");
    gpmc_send('1',x"2D38",x"2D00");
    gpmc_send('1',x"2D39",x"0012");
    gpmc_send('1',x"2D3A",x"2E00");
    gpmc_send('1',x"2D3B",x"0011");
    gpmc_send('1',x"2D3C",x"2F00");
    gpmc_send('1',x"2D3D",x"0010");
    gpmc_send('1',x"2D3E",x"3000");
    gpmc_send('1',x"2D3F",x"000F");
    gpmc_send('1',x"2D40",x"3100");
    gpmc_send('1',x"2D41",x"000E");
    gpmc_send('1',x"2D42",x"3200");
    gpmc_send('1',x"2D43",x"000D");
    gpmc_send('1',x"2D44",x"3300");
    gpmc_send('1',x"2D45",x"000C");
    gpmc_send('1',x"2D46",x"3400");
    gpmc_send('1',x"2D47",x"000B");
    gpmc_send('1',x"2D48",x"3500");
    gpmc_send('1',x"2D49",x"000A");
    gpmc_send('1',x"2D4A",x"3600");
    gpmc_send('1',x"2D4B",x"0009");
    gpmc_send('1',x"2D4C",x"3700");
    gpmc_send('1',x"2D4D",x"0008");
    gpmc_send('1',x"2D4E",x"3800");
    gpmc_send('1',x"2D4F",x"0007");
    gpmc_send('1',x"2D50",x"3900");
    gpmc_send('1',x"2D51",x"0006");
    gpmc_send('1',x"2D52",x"3A00");
    gpmc_send('1',x"2D53",x"0005");
    gpmc_send('1',x"2D54",x"3B00");
    gpmc_send('1',x"2D55",x"0004");
    gpmc_send('1',x"2D56",x"3C00");
    gpmc_send('1',x"2D57",x"0003");
    gpmc_send('1',x"2D58",x"3D00");
    gpmc_send('1',x"2D59",x"0002");
    gpmc_send('1',x"2D5A",x"3E00");
    gpmc_send('1',x"2D5B",x"0001");
    gpmc_send('1',x"2D5C",x"3F00");
    gpmc_send('1',x"2D5D",x"0000");
    gpmc_send('1',x"2D5E",x"3F01");
    gpmc_send('1',x"2D5F",x"0000");
    gpmc_send('1',x"2D60",x"3E02");
    gpmc_send('1',x"2D61",x"0000");
    gpmc_send('1',x"2D62",x"3D03");
    gpmc_send('1',x"2D63",x"0000");
    gpmc_send('1',x"2D64",x"3C04");
    gpmc_send('1',x"2D65",x"0000");
    gpmc_send('1',x"2D66",x"3B05");
    gpmc_send('1',x"2D67",x"0000");
    gpmc_send('1',x"2D68",x"3A06");
    gpmc_send('1',x"2D69",x"0000");
    gpmc_send('1',x"2D6A",x"3907");
    gpmc_send('1',x"2D6B",x"0000");
    gpmc_send('1',x"2D6C",x"3808");
    gpmc_send('1',x"2D6D",x"0000");
    gpmc_send('1',x"2D6E",x"3709");
    gpmc_send('1',x"2D6F",x"0000");
    gpmc_send('1',x"2D70",x"360A");
    gpmc_send('1',x"2D71",x"0000");
    gpmc_send('1',x"2D72",x"350B");
    gpmc_send('1',x"2D73",x"0000");
    gpmc_send('1',x"2D74",x"340C");
    gpmc_send('1',x"2D75",x"0000");
    gpmc_send('1',x"2D76",x"330D");
    gpmc_send('1',x"2D77",x"0000");
    gpmc_send('1',x"2D78",x"320E");
    gpmc_send('1',x"2D79",x"0000");
    gpmc_send('1',x"2D7A",x"310F");
    gpmc_send('1',x"2D7B",x"0000");
    gpmc_send('1',x"2D7C",x"3010");
    gpmc_send('1',x"2D7D",x"0000");
    gpmc_send('1',x"2D7E",x"2F11");
    gpmc_send('1',x"2D7F",x"0000");
    gpmc_send('1',x"2D80",x"2E12");
    gpmc_send('1',x"2D81",x"0000");
    gpmc_send('1',x"2D82",x"2D13");
    gpmc_send('1',x"2D83",x"0000");
    gpmc_send('1',x"2D84",x"2C14");
    gpmc_send('1',x"2D85",x"0000");
    gpmc_send('1',x"2D86",x"2B15");
    gpmc_send('1',x"2D87",x"0000");
    gpmc_send('1',x"2D88",x"2A16");
    gpmc_send('1',x"2D89",x"0000");
    gpmc_send('1',x"2D8A",x"2917");
    gpmc_send('1',x"2D8B",x"0000");
    gpmc_send('1',x"2D8C",x"2818");
    gpmc_send('1',x"2D8D",x"0000");
    gpmc_send('1',x"2D8E",x"2719");
    gpmc_send('1',x"2D8F",x"0000");
    gpmc_send('1',x"2D90",x"261A");
    gpmc_send('1',x"2D91",x"0000");
    gpmc_send('1',x"2D92",x"251B");
    gpmc_send('1',x"2D93",x"0000");
    gpmc_send('1',x"2D94",x"241C");
    gpmc_send('1',x"2D95",x"0000");
    gpmc_send('1',x"2D96",x"231D");
    gpmc_send('1',x"2D97",x"0000");
    gpmc_send('1',x"2D98",x"221E");
    gpmc_send('1',x"2D99",x"0000");
    gpmc_send('1',x"2D9A",x"211F");
    gpmc_send('1',x"2D9B",x"0000");
    gpmc_send('1',x"2D9C",x"2020");
    gpmc_send('1',x"2D9D",x"0000");
    gpmc_send('1',x"2D9E",x"1F21");
    gpmc_send('1',x"2D9F",x"0000");
    gpmc_send('1',x"2DA0",x"1E22");
    gpmc_send('1',x"2DA1",x"0000");
    gpmc_send('1',x"2DA2",x"1D23");
    gpmc_send('1',x"2DA3",x"0000");
    gpmc_send('1',x"2DA4",x"1C24");
    gpmc_send('1',x"2DA5",x"0000");
    gpmc_send('1',x"2DA6",x"1B25");
    gpmc_send('1',x"2DA7",x"0000");
    gpmc_send('1',x"2DA8",x"1A26");
    gpmc_send('1',x"2DA9",x"0000");
    gpmc_send('1',x"2DAA",x"1927");
    gpmc_send('1',x"2DAB",x"0000");
    gpmc_send('1',x"2DAC",x"1828");
    gpmc_send('1',x"2DAD",x"0000");
    gpmc_send('1',x"2DAE",x"1729");
    gpmc_send('1',x"2DAF",x"0000");
    gpmc_send('1',x"2DB0",x"162A");
    gpmc_send('1',x"2DB1",x"0000");
    gpmc_send('1',x"2DB2",x"152B");
    gpmc_send('1',x"2DB3",x"0000");
    gpmc_send('1',x"2DB4",x"142C");
    gpmc_send('1',x"2DB5",x"0000");
    gpmc_send('1',x"2DB6",x"132D");
    gpmc_send('1',x"2DB7",x"0000");
    gpmc_send('1',x"2DB8",x"122E");
    gpmc_send('1',x"2DB9",x"0000");
    gpmc_send('1',x"2DBA",x"112F");
    gpmc_send('1',x"2DBB",x"0000");
    gpmc_send('1',x"2DBC",x"1030");
    gpmc_send('1',x"2DBD",x"0000");
    gpmc_send('1',x"2DBE",x"0F31");
    gpmc_send('1',x"2DBF",x"0000");
    gpmc_send('1',x"2DC0",x"0E32");
    gpmc_send('1',x"2DC1",x"0000");
    gpmc_send('1',x"2DC2",x"0D33");
    gpmc_send('1',x"2DC3",x"0000");
    gpmc_send('1',x"2DC4",x"0C34");
    gpmc_send('1',x"2DC5",x"0000");
    gpmc_send('1',x"2DC6",x"0B35");
    gpmc_send('1',x"2DC7",x"0000");
    gpmc_send('1',x"2DC8",x"0A36");
    gpmc_send('1',x"2DC9",x"0000");
    gpmc_send('1',x"2DCA",x"0937");
    gpmc_send('1',x"2DCB",x"0000");
    gpmc_send('1',x"2DCC",x"0838");
    gpmc_send('1',x"2DCD",x"0000");
    gpmc_send('1',x"2DCE",x"0739");
    gpmc_send('1',x"2DCF",x"0000");
    gpmc_send('1',x"2DD0",x"063A");
    gpmc_send('1',x"2DD1",x"0000");
    gpmc_send('1',x"2DD2",x"053B");
    gpmc_send('1',x"2DD3",x"0000");
    gpmc_send('1',x"2DD4",x"043C");
    gpmc_send('1',x"2DD5",x"0000");
    gpmc_send('1',x"2DD6",x"033D");
    gpmc_send('1',x"2DD7",x"0000");
    gpmc_send('1',x"2DD8",x"023E");
    gpmc_send('1',x"2DD9",x"0000");
    gpmc_send('1',x"2DDA",x"013F");
    gpmc_send('1',x"2DDB",x"0000");
    gpmc_send('1',x"2DDC",x"003F");
    gpmc_send('1',x"2DDD",x"0000");
    gpmc_send('1',x"2DDE",x"003E");
    gpmc_send('1',x"2DDF",x"0001");
    gpmc_send('1',x"2DE0",x"003D");
    gpmc_send('1',x"2DE1",x"0002");
    gpmc_send('1',x"2DE2",x"003C");
    gpmc_send('1',x"2DE3",x"0003");
    gpmc_send('1',x"2DE4",x"003B");
    gpmc_send('1',x"2DE5",x"0004");
    gpmc_send('1',x"2DE6",x"003A");
    gpmc_send('1',x"2DE7",x"0005");
    gpmc_send('1',x"2DE8",x"0039");
    gpmc_send('1',x"2DE9",x"0006");
    gpmc_send('1',x"2DEA",x"0038");
    gpmc_send('1',x"2DEB",x"0007");
    gpmc_send('1',x"2DEC",x"0037");
    gpmc_send('1',x"2DED",x"0008");
    gpmc_send('1',x"2DEE",x"0036");
    gpmc_send('1',x"2DEF",x"0009");
    gpmc_send('1',x"2DF0",x"0035");
    gpmc_send('1',x"2DF1",x"000A");
    gpmc_send('1',x"2DF2",x"0034");
    gpmc_send('1',x"2DF3",x"000B");
    gpmc_send('1',x"2DF4",x"0033");
    gpmc_send('1',x"2DF5",x"000C");
    gpmc_send('1',x"2DF6",x"0032");
    gpmc_send('1',x"2DF7",x"000D");
    gpmc_send('1',x"2DF8",x"0031");
    gpmc_send('1',x"2DF9",x"000E");
    gpmc_send('1',x"2DFA",x"0030");
    gpmc_send('1',x"2DFB",x"000F");
    gpmc_send('1',x"2DFC",x"002F");
    gpmc_send('1',x"2DFD",x"0010");
    gpmc_send('1',x"2DFE",x"002E");
    gpmc_send('1',x"2DFF",x"0011");
    gpmc_send('1',x"2E00",x"002D");
    gpmc_send('1',x"2E01",x"0012");
    gpmc_send('1',x"2E02",x"002C");
    gpmc_send('1',x"2E03",x"0013");
    gpmc_send('1',x"2E04",x"002B");
    gpmc_send('1',x"2E05",x"0014");
    gpmc_send('1',x"2E06",x"002A");
    gpmc_send('1',x"2E07",x"0015");
    gpmc_send('1',x"2E08",x"0029");
    gpmc_send('1',x"2E09",x"0016");
    gpmc_send('1',x"2E0A",x"0028");
    gpmc_send('1',x"2E0B",x"0017");
    gpmc_send('1',x"2E0C",x"0027");
    gpmc_send('1',x"2E0D",x"0018");
    gpmc_send('1',x"2E0E",x"0026");
    gpmc_send('1',x"2E0F",x"0019");
    gpmc_send('1',x"2E10",x"0025");
    gpmc_send('1',x"2E11",x"001A");
    gpmc_send('1',x"2E12",x"0024");
    gpmc_send('1',x"2E13",x"001B");
    gpmc_send('1',x"2E14",x"0023");
    gpmc_send('1',x"2E15",x"001C");
    gpmc_send('1',x"2E16",x"0022");
    gpmc_send('1',x"2E17",x"001D");
    gpmc_send('1',x"2E18",x"0021");
    gpmc_send('1',x"2E19",x"001E");
    gpmc_send('1',x"2E1A",x"0020");
    gpmc_send('1',x"2E1B",x"001F");
    gpmc_send('1',x"2E1C",x"001F");
    gpmc_send('1',x"2E1D",x"0020");
    gpmc_send('1',x"2E1E",x"001E");
    gpmc_send('1',x"2E1F",x"0021");
    gpmc_send('1',x"2E20",x"001D");
    gpmc_send('1',x"2E21",x"0022");
    gpmc_send('1',x"2E22",x"001C");
    gpmc_send('1',x"2E23",x"0023");
    gpmc_send('1',x"2E24",x"001B");
    gpmc_send('1',x"2E25",x"0024");
    gpmc_send('1',x"2E26",x"001A");
    gpmc_send('1',x"2E27",x"0025");
    gpmc_send('1',x"2E28",x"0019");
    gpmc_send('1',x"2E29",x"0026");
    gpmc_send('1',x"2E2A",x"0018");
    gpmc_send('1',x"2E2B",x"0027");
    gpmc_send('1',x"2E2C",x"0017");
    gpmc_send('1',x"2E2D",x"0028");
    gpmc_send('1',x"2E2E",x"0016");
    gpmc_send('1',x"2E2F",x"0029");
    gpmc_send('1',x"2E30",x"0015");
    gpmc_send('1',x"2E31",x"002A");
    gpmc_send('1',x"2E32",x"0014");
    gpmc_send('1',x"2E33",x"002B");
    gpmc_send('1',x"2E34",x"0013");
    gpmc_send('1',x"2E35",x"002C");
    gpmc_send('1',x"2E36",x"0012");
    gpmc_send('1',x"2E37",x"002D");
    gpmc_send('1',x"2E38",x"0011");
    gpmc_send('1',x"2E39",x"002E");
    gpmc_send('1',x"2E3A",x"0010");
    gpmc_send('1',x"2E3B",x"002F");
    gpmc_send('1',x"2E3C",x"000F");
    gpmc_send('1',x"2E3D",x"0030");
    gpmc_send('1',x"2E3E",x"000E");
    gpmc_send('1',x"2E3F",x"0031");
    gpmc_send('1',x"2E40",x"000D");
    gpmc_send('1',x"2E41",x"0032");
    gpmc_send('1',x"2E42",x"000C");
    gpmc_send('1',x"2E43",x"0033");
    gpmc_send('1',x"2E44",x"000B");
    gpmc_send('1',x"2E45",x"0034");
    gpmc_send('1',x"2E46",x"000A");
    gpmc_send('1',x"2E47",x"0035");
    gpmc_send('1',x"2E48",x"0009");
    gpmc_send('1',x"2E49",x"0036");
    gpmc_send('1',x"2E4A",x"0008");
    gpmc_send('1',x"2E4B",x"0037");
    gpmc_send('1',x"2E4C",x"0007");
    gpmc_send('1',x"2E4D",x"0038");
    gpmc_send('1',x"2E4E",x"0006");
    gpmc_send('1',x"2E4F",x"0039");
    gpmc_send('1',x"2E50",x"0005");
    gpmc_send('1',x"2E51",x"003A");
    gpmc_send('1',x"2E52",x"0004");
    gpmc_send('1',x"2E53",x"003B");
    gpmc_send('1',x"2E54",x"0003");
    gpmc_send('1',x"2E55",x"003C");
    gpmc_send('1',x"2E56",x"0002");
    gpmc_send('1',x"2E57",x"003D");
    gpmc_send('1',x"2E58",x"0001");
    gpmc_send('1',x"2E59",x"003E");
    gpmc_send('1',x"2E5A",x"0000");
    gpmc_send('1',x"2E5B",x"003F");
    gpmc_send('1',x"2E5C",x"0100");
    gpmc_send('1',x"2E5D",x"003E");
    gpmc_send('1',x"2E5E",x"0200");
    gpmc_send('1',x"2E5F",x"003D");
    gpmc_send('1',x"2E60",x"0300");
    gpmc_send('1',x"2E61",x"003C");
    gpmc_send('1',x"2E62",x"0400");
    gpmc_send('1',x"2E63",x"003B");
    gpmc_send('1',x"2E64",x"0500");
    gpmc_send('1',x"2E65",x"003A");
    gpmc_send('1',x"2E66",x"0600");
    gpmc_send('1',x"2E67",x"0039");
    gpmc_send('1',x"2E68",x"0700");
    gpmc_send('1',x"2E69",x"0038");
    gpmc_send('1',x"2E6A",x"0800");
    gpmc_send('1',x"2E6B",x"0037");
    gpmc_send('1',x"2E6C",x"0900");
    gpmc_send('1',x"2E6D",x"0036");
    gpmc_send('1',x"2E6E",x"0A00");
    gpmc_send('1',x"2E6F",x"0035");
    gpmc_send('1',x"2E70",x"0B00");
    gpmc_send('1',x"2E71",x"0034");
    gpmc_send('1',x"2E72",x"0C00");
    gpmc_send('1',x"2E73",x"0033");
    gpmc_send('1',x"2E74",x"0D00");
    gpmc_send('1',x"2E75",x"0032");
    gpmc_send('1',x"2E76",x"0E00");
    gpmc_send('1',x"2E77",x"0031");
    gpmc_send('1',x"2E78",x"0F00");
    gpmc_send('1',x"2E79",x"0030");
    gpmc_send('1',x"2E7A",x"1000");
    gpmc_send('1',x"2E7B",x"002F");
    gpmc_send('1',x"2E7C",x"1100");
    gpmc_send('1',x"2E7D",x"002E");
    gpmc_send('1',x"2E7E",x"1200");
    gpmc_send('1',x"2E7F",x"002D");
    gpmc_send('1',x"2E80",x"1300");
    gpmc_send('1',x"2E81",x"002C");
    gpmc_send('1',x"2E82",x"1400");
    gpmc_send('1',x"2E83",x"002B");
    gpmc_send('1',x"2E84",x"1500");
    gpmc_send('1',x"2E85",x"002A");
    gpmc_send('1',x"2E86",x"1600");
    gpmc_send('1',x"2E87",x"0029");
    gpmc_send('1',x"2E88",x"1700");
    gpmc_send('1',x"2E89",x"0028");
    gpmc_send('1',x"2E8A",x"1800");
    gpmc_send('1',x"2E8B",x"0027");
    gpmc_send('1',x"2E8C",x"1900");
    gpmc_send('1',x"2E8D",x"0026");
    gpmc_send('1',x"2E8E",x"1A00");
    gpmc_send('1',x"2E8F",x"0025");
    gpmc_send('1',x"2E90",x"1B00");
    gpmc_send('1',x"2E91",x"0024");
    gpmc_send('1',x"2E92",x"1C00");
    gpmc_send('1',x"2E93",x"0023");
    gpmc_send('1',x"2E94",x"1D00");
    gpmc_send('1',x"2E95",x"0022");
    gpmc_send('1',x"2E96",x"1E00");
    gpmc_send('1',x"2E97",x"0021");
    gpmc_send('1',x"2E98",x"1F00");
    gpmc_send('1',x"2E99",x"0020");
    gpmc_send('1',x"2E9A",x"2000");
    gpmc_send('1',x"2E9B",x"001F");
    gpmc_send('1',x"2E9C",x"2100");
    gpmc_send('1',x"2E9D",x"001E");
    gpmc_send('1',x"2E9E",x"2200");
    gpmc_send('1',x"2E9F",x"001D");
    gpmc_send('1',x"2EA0",x"2300");
    gpmc_send('1',x"2EA1",x"001C");
    gpmc_send('1',x"2EA2",x"2400");
    gpmc_send('1',x"2EA3",x"001B");
    gpmc_send('1',x"2EA4",x"2500");
    gpmc_send('1',x"2EA5",x"001A");
    gpmc_send('1',x"2EA6",x"2600");
    gpmc_send('1',x"2EA7",x"0019");
    gpmc_send('1',x"2EA8",x"2700");
    gpmc_send('1',x"2EA9",x"0018");
    gpmc_send('1',x"2EAA",x"2800");
    gpmc_send('1',x"2EAB",x"0017");
    gpmc_send('1',x"2EAC",x"2900");
    gpmc_send('1',x"2EAD",x"0016");
    gpmc_send('1',x"2EAE",x"2A00");
    gpmc_send('1',x"2EAF",x"0015");
    gpmc_send('1',x"2EB0",x"2B00");
    gpmc_send('1',x"2EB1",x"0014");
    gpmc_send('1',x"2EB2",x"2C00");
    gpmc_send('1',x"2EB3",x"0013");
    gpmc_send('1',x"2EB4",x"2D00");
    gpmc_send('1',x"2EB5",x"0012");
    gpmc_send('1',x"2EB6",x"2E00");
    gpmc_send('1',x"2EB7",x"0011");
    gpmc_send('1',x"2EB8",x"2F00");
    gpmc_send('1',x"2EB9",x"0010");
    gpmc_send('1',x"2EBA",x"3000");
    gpmc_send('1',x"2EBB",x"000F");
    gpmc_send('1',x"2EBC",x"3100");
    gpmc_send('1',x"2EBD",x"000E");
    gpmc_send('1',x"2EBE",x"3200");
    gpmc_send('1',x"2EBF",x"000D");
    gpmc_send('1',x"2EC0",x"3300");
    gpmc_send('1',x"2EC1",x"000C");
    gpmc_send('1',x"2EC2",x"3400");
    gpmc_send('1',x"2EC3",x"000B");
    gpmc_send('1',x"2EC4",x"3500");
    gpmc_send('1',x"2EC5",x"000A");
    gpmc_send('1',x"2EC6",x"3600");
    gpmc_send('1',x"2EC7",x"0009");
    gpmc_send('1',x"2EC8",x"3700");
    gpmc_send('1',x"2EC9",x"0008");
    gpmc_send('1',x"2ECA",x"3800");
    gpmc_send('1',x"2ECB",x"0007");
    gpmc_send('1',x"2ECC",x"3900");
    gpmc_send('1',x"2ECD",x"0006");
    gpmc_send('1',x"2ECE",x"3A00");
    gpmc_send('1',x"2ECF",x"0005");
    gpmc_send('1',x"2ED0",x"3B00");
    gpmc_send('1',x"2ED1",x"0004");
    gpmc_send('1',x"2ED2",x"3C00");
    gpmc_send('1',x"2ED3",x"0003");
    gpmc_send('1',x"2ED4",x"3D00");
    gpmc_send('1',x"2ED5",x"0002");
    gpmc_send('1',x"2ED6",x"3E00");
    gpmc_send('1',x"2ED7",x"0001");
    gpmc_send('1',x"2ED8",x"3F00");
    gpmc_send('1',x"2ED9",x"0000");
    gpmc_send('1',x"2EDA",x"3F01");
    gpmc_send('1',x"2EDB",x"0000");
    gpmc_send('1',x"2EDC",x"3E02");
    gpmc_send('1',x"2EDD",x"0000");
    gpmc_send('1',x"2EDE",x"3D03");
    gpmc_send('1',x"2EDF",x"0000");
    gpmc_send('1',x"2EE0",x"3C04");
    gpmc_send('1',x"2EE1",x"0000");
    gpmc_send('1',x"2EE2",x"3B05");
    gpmc_send('1',x"2EE3",x"0000");
    gpmc_send('1',x"2EE4",x"3A06");
    gpmc_send('1',x"2EE5",x"0000");
    gpmc_send('1',x"2EE6",x"3907");
    gpmc_send('1',x"2EE7",x"0000");
    gpmc_send('1',x"2EE8",x"3808");
    gpmc_send('1',x"2EE9",x"0000");
    gpmc_send('1',x"2EEA",x"3709");
    gpmc_send('1',x"2EEB",x"0000");
    gpmc_send('1',x"2EEC",x"360A");
    gpmc_send('1',x"2EED",x"0000");
    gpmc_send('1',x"2EEE",x"350B");
    gpmc_send('1',x"2EEF",x"0000");
    gpmc_send('1',x"2EF0",x"340C");
    gpmc_send('1',x"2EF1",x"0000");
    gpmc_send('1',x"2EF2",x"330D");
    gpmc_send('1',x"2EF3",x"0000");
    gpmc_send('1',x"2EF4",x"320E");
    gpmc_send('1',x"2EF5",x"0000");
    gpmc_send('1',x"2EF6",x"310F");
    gpmc_send('1',x"2EF7",x"0000");
    gpmc_send('1',x"2EF8",x"3010");
    gpmc_send('1',x"2EF9",x"0000");
    gpmc_send('1',x"2EFA",x"2F11");
    gpmc_send('1',x"2EFB",x"0000");
    gpmc_send('1',x"2EFC",x"2E12");
    gpmc_send('1',x"2EFD",x"0000");
    gpmc_send('1',x"2EFE",x"2D13");
    gpmc_send('1',x"2EFF",x"0000");
    gpmc_send('1',x"2F00",x"2C14");
    gpmc_send('1',x"2F01",x"0000");
    gpmc_send('1',x"2F02",x"2B15");
    gpmc_send('1',x"2F03",x"0000");
    gpmc_send('1',x"2F04",x"2A16");
    gpmc_send('1',x"2F05",x"0000");
    gpmc_send('1',x"2F06",x"2917");
    gpmc_send('1',x"2F07",x"0000");
    gpmc_send('1',x"2F08",x"2818");
    gpmc_send('1',x"2F09",x"0000");
    gpmc_send('1',x"2F0A",x"2719");
    gpmc_send('1',x"2F0B",x"0000");
    gpmc_send('1',x"2F0C",x"261A");
    gpmc_send('1',x"2F0D",x"0000");
    gpmc_send('1',x"2F0E",x"251B");
    gpmc_send('1',x"2F0F",x"0000");
    gpmc_send('1',x"2F10",x"241C");
    gpmc_send('1',x"2F11",x"0000");
    gpmc_send('1',x"2F12",x"231D");
    gpmc_send('1',x"2F13",x"0000");
    gpmc_send('1',x"2F14",x"221E");
    gpmc_send('1',x"2F15",x"0000");
    gpmc_send('1',x"2F16",x"211F");
    gpmc_send('1',x"2F17",x"0000");
    gpmc_send('1',x"2F18",x"2020");
    gpmc_send('1',x"2F19",x"0000");
    gpmc_send('1',x"2F1A",x"1F21");
    gpmc_send('1',x"2F1B",x"0000");
    gpmc_send('1',x"2F1C",x"1E22");
    gpmc_send('1',x"2F1D",x"0000");
    gpmc_send('1',x"2F1E",x"1D23");
    gpmc_send('1',x"2F1F",x"0000");
    gpmc_send('1',x"2F20",x"1C24");
    gpmc_send('1',x"2F21",x"0000");
    gpmc_send('1',x"2F22",x"1B25");
    gpmc_send('1',x"2F23",x"0000");
    gpmc_send('1',x"2F24",x"1A26");
    gpmc_send('1',x"2F25",x"0000");
    gpmc_send('1',x"2F26",x"1927");
    gpmc_send('1',x"2F27",x"0000");
    gpmc_send('1',x"2F28",x"1828");
    gpmc_send('1',x"2F29",x"0000");
    gpmc_send('1',x"2F2A",x"1729");
    gpmc_send('1',x"2F2B",x"0000");
    gpmc_send('1',x"2F2C",x"162A");
    gpmc_send('1',x"2F2D",x"0000");
    gpmc_send('1',x"2F2E",x"152B");
    gpmc_send('1',x"2F2F",x"0000");
    gpmc_send('1',x"2F30",x"142C");
    gpmc_send('1',x"2F31",x"0000");
    gpmc_send('1',x"2F32",x"132D");
    gpmc_send('1',x"2F33",x"0000");
    gpmc_send('1',x"2F34",x"122E");
    gpmc_send('1',x"2F35",x"0000");
    gpmc_send('1',x"2F36",x"112F");
    gpmc_send('1',x"2F37",x"0000");
    gpmc_send('1',x"2F38",x"1030");
    gpmc_send('1',x"2F39",x"0000");
    gpmc_send('1',x"2F3A",x"0F31");
    gpmc_send('1',x"2F3B",x"0000");
    gpmc_send('1',x"2F3C",x"0E32");
    gpmc_send('1',x"2F3D",x"0000");
    gpmc_send('1',x"2F3E",x"0D33");
    gpmc_send('1',x"2F3F",x"0000");
    gpmc_send('1',x"2F40",x"0C34");
    gpmc_send('1',x"2F41",x"0000");
    gpmc_send('1',x"2F42",x"0B35");
    gpmc_send('1',x"2F43",x"0000");
    gpmc_send('1',x"2F44",x"0A36");
    gpmc_send('1',x"2F45",x"0000");
    gpmc_send('1',x"2F46",x"0937");
    gpmc_send('1',x"2F47",x"0000");
    gpmc_send('1',x"2F48",x"0838");
    gpmc_send('1',x"2F49",x"0000");
    gpmc_send('1',x"2F4A",x"0739");
    gpmc_send('1',x"2F4B",x"0000");
    gpmc_send('1',x"2F4C",x"063A");
    gpmc_send('1',x"2F4D",x"0000");
    gpmc_send('1',x"2F4E",x"053B");
    gpmc_send('1',x"2F4F",x"0000");
    gpmc_send('1',x"2F50",x"043C");
    gpmc_send('1',x"2F51",x"0000");
    gpmc_send('1',x"2F52",x"033D");
    gpmc_send('1',x"2F53",x"0000");
    gpmc_send('1',x"2F54",x"023E");
    gpmc_send('1',x"2F55",x"0000");
    gpmc_send('1',x"2F56",x"013F");
    gpmc_send('1',x"2F57",x"0000");
    gpmc_send('1',x"2F58",x"003F");
    gpmc_send('1',x"2F59",x"0000");
    gpmc_send('1',x"2F5A",x"003E");
    gpmc_send('1',x"2F5B",x"0001");
    gpmc_send('1',x"2F5C",x"003D");
    gpmc_send('1',x"2F5D",x"0002");
    gpmc_send('1',x"2F5E",x"003C");
    gpmc_send('1',x"2F5F",x"0003");
    gpmc_send('1',x"2F60",x"003B");
    gpmc_send('1',x"2F61",x"0004");
    gpmc_send('1',x"2F62",x"003A");
    gpmc_send('1',x"2F63",x"0005");
    gpmc_send('1',x"2F64",x"0039");
    gpmc_send('1',x"2F65",x"0006");
    gpmc_send('1',x"2F66",x"0038");
    gpmc_send('1',x"2F67",x"0007");
    gpmc_send('1',x"2F68",x"0037");
    gpmc_send('1',x"2F69",x"0008");
    gpmc_send('1',x"2F6A",x"0036");
    gpmc_send('1',x"2F6B",x"0009");
    gpmc_send('1',x"2F6C",x"0035");
    gpmc_send('1',x"2F6D",x"000A");
    gpmc_send('1',x"2F6E",x"0034");
    gpmc_send('1',x"2F6F",x"000B");
    gpmc_send('1',x"2F70",x"0033");
    gpmc_send('1',x"2F71",x"000C");
    gpmc_send('1',x"2F72",x"0032");
    gpmc_send('1',x"2F73",x"000D");
    gpmc_send('1',x"2F74",x"0031");
    gpmc_send('1',x"2F75",x"000E");
    gpmc_send('1',x"2F76",x"0030");
    gpmc_send('1',x"2F77",x"000F");
    gpmc_send('1',x"2F78",x"002F");
    gpmc_send('1',x"2F79",x"0010");
    gpmc_send('1',x"2F7A",x"002E");
    gpmc_send('1',x"2F7B",x"0011");
    gpmc_send('1',x"2F7C",x"002D");
    gpmc_send('1',x"2F7D",x"0012");
    gpmc_send('1',x"2F7E",x"002C");
    gpmc_send('1',x"2F7F",x"0013");
    gpmc_send('1',x"2F80",x"002B");
    gpmc_send('1',x"2F81",x"0014");
    gpmc_send('1',x"2F82",x"002A");
    gpmc_send('1',x"2F83",x"0015");
    gpmc_send('1',x"2F84",x"0029");
    gpmc_send('1',x"2F85",x"0016");
    gpmc_send('1',x"2F86",x"0028");
    gpmc_send('1',x"2F87",x"0017");
    gpmc_send('1',x"2F88",x"0027");
    gpmc_send('1',x"2F89",x"0018");
    gpmc_send('1',x"2F8A",x"0026");
    gpmc_send('1',x"2F8B",x"0019");
    gpmc_send('1',x"2F8C",x"0025");
    gpmc_send('1',x"2F8D",x"001A");
    gpmc_send('1',x"2F8E",x"0024");
    gpmc_send('1',x"2F8F",x"001B");
    gpmc_send('1',x"2F90",x"0023");
    gpmc_send('1',x"2F91",x"001C");
    gpmc_send('1',x"2F92",x"0022");
    gpmc_send('1',x"2F93",x"001D");
    gpmc_send('1',x"2F94",x"0021");
    gpmc_send('1',x"2F95",x"001E");
    gpmc_send('1',x"2F96",x"0020");
    gpmc_send('1',x"2F97",x"001F");
    gpmc_send('1',x"2F98",x"001F");
    gpmc_send('1',x"2F99",x"0020");
    gpmc_send('1',x"2F9A",x"001E");
    gpmc_send('1',x"2F9B",x"0021");
    gpmc_send('1',x"2F9C",x"001D");
    gpmc_send('1',x"2F9D",x"0022");
    gpmc_send('1',x"2F9E",x"001C");
    gpmc_send('1',x"2F9F",x"0023");
    gpmc_send('1',x"2FA0",x"001B");
    gpmc_send('1',x"2FA1",x"0024");
    gpmc_send('1',x"2FA2",x"001A");
    gpmc_send('1',x"2FA3",x"0025");
    gpmc_send('1',x"2FA4",x"0019");
    gpmc_send('1',x"2FA5",x"0026");
    gpmc_send('1',x"2FA6",x"0018");
    gpmc_send('1',x"2FA7",x"0027");
    gpmc_send('1',x"2FA8",x"0017");
    gpmc_send('1',x"2FA9",x"0028");
    gpmc_send('1',x"2FAA",x"0016");
    gpmc_send('1',x"2FAB",x"0029");
    gpmc_send('1',x"2FAC",x"0015");
    gpmc_send('1',x"2FAD",x"002A");
    gpmc_send('1',x"2FAE",x"0014");
    gpmc_send('1',x"2FAF",x"002B");
    gpmc_send('1',x"2FB0",x"0013");
    gpmc_send('1',x"2FB1",x"002C");
    gpmc_send('1',x"2FB2",x"0012");
    gpmc_send('1',x"2FB3",x"002D");
    gpmc_send('1',x"2FB4",x"0011");
    gpmc_send('1',x"2FB5",x"002E");
    gpmc_send('1',x"2FB6",x"0010");
    gpmc_send('1',x"2FB7",x"002F");
    gpmc_send('1',x"2FB8",x"000F");
    gpmc_send('1',x"2FB9",x"0030");
    gpmc_send('1',x"2FBA",x"000E");
    gpmc_send('1',x"2FBB",x"0031");
    gpmc_send('1',x"2FBC",x"000D");
    gpmc_send('1',x"2FBD",x"0032");
    gpmc_send('1',x"2FBE",x"000C");
    gpmc_send('1',x"2FBF",x"0033");
    gpmc_send('1',x"2FC0",x"000B");
    gpmc_send('1',x"2FC1",x"0034");
    gpmc_send('1',x"2FC2",x"000A");
    gpmc_send('1',x"2FC3",x"0035");
    gpmc_send('1',x"2FC4",x"0009");
    gpmc_send('1',x"2FC5",x"0036");
    gpmc_send('1',x"2FC6",x"0008");
    gpmc_send('1',x"2FC7",x"0037");
    gpmc_send('1',x"2FC8",x"0007");
    gpmc_send('1',x"2FC9",x"0038");
    gpmc_send('1',x"2FCA",x"0006");
    gpmc_send('1',x"2FCB",x"0039");
    gpmc_send('1',x"2FCC",x"0005");
    gpmc_send('1',x"2FCD",x"003A");
    gpmc_send('1',x"2FCE",x"0004");
    gpmc_send('1',x"2FCF",x"003B");
    gpmc_send('1',x"2FD0",x"0003");
    gpmc_send('1',x"2FD1",x"003C");
    gpmc_send('1',x"2FD2",x"0002");
    gpmc_send('1',x"2FD3",x"003D");
    gpmc_send('1',x"2FD4",x"0001");
    gpmc_send('1',x"2FD5",x"003E");
    gpmc_send('1',x"2FD6",x"0000");
    gpmc_send('1',x"2FD7",x"003F");
    gpmc_send('1',x"2FD8",x"0100");
    gpmc_send('1',x"2FD9",x"003E");
    gpmc_send('1',x"2FDA",x"0200");
    gpmc_send('1',x"2FDB",x"003D");
    gpmc_send('1',x"2FDC",x"0300");
    gpmc_send('1',x"2FDD",x"003C");
    gpmc_send('1',x"2FDE",x"0400");
    gpmc_send('1',x"2FDF",x"003B");
    gpmc_send('1',x"2FE0",x"0500");
    gpmc_send('1',x"2FE1",x"003A");
    gpmc_send('1',x"2FE2",x"0600");
    gpmc_send('1',x"2FE3",x"0039");
    gpmc_send('1',x"2FE4",x"0700");
    gpmc_send('1',x"2FE5",x"0038");
    gpmc_send('1',x"2FE6",x"0800");
    gpmc_send('1',x"2FE7",x"0037");
    gpmc_send('1',x"2FE8",x"0900");
    gpmc_send('1',x"2FE9",x"0036");
    gpmc_send('1',x"2FEA",x"0A00");
    gpmc_send('1',x"2FEB",x"0035");
    gpmc_send('1',x"2FEC",x"0B00");
    gpmc_send('1',x"2FED",x"0034");
    gpmc_send('1',x"2FEE",x"0C00");
    gpmc_send('1',x"2FEF",x"0033");
    gpmc_send('1',x"2FF0",x"0D00");
    gpmc_send('1',x"2FF1",x"0032");
    gpmc_send('1',x"2FF2",x"0E00");
    gpmc_send('1',x"2FF3",x"0031");
    gpmc_send('1',x"2FF4",x"0F00");
    gpmc_send('1',x"2FF5",x"0030");
    gpmc_send('1',x"2FF6",x"1000");
    gpmc_send('1',x"2FF7",x"002F");
    gpmc_send('1',x"2FF8",x"1100");
    gpmc_send('1',x"2FF9",x"002E");
    gpmc_send('1',x"2FFA",x"1200");
    gpmc_send('1',x"2FFB",x"002D");
    gpmc_send('1',x"2FFC",x"1300");
    gpmc_send('1',x"2FFD",x"002C");
    gpmc_send('1',x"2FFE",x"1400");
    gpmc_send('1',x"2FFF",x"002B");
    gpmc_send('1',x"3000",x"1500");
    gpmc_send('1',x"3001",x"002A");
    gpmc_send('1',x"3002",x"1600");
    gpmc_send('1',x"3003",x"0029");
    gpmc_send('1',x"3004",x"1700");
    gpmc_send('1',x"3005",x"0028");
    gpmc_send('1',x"3006",x"1800");
    gpmc_send('1',x"3007",x"0027");
    gpmc_send('1',x"3008",x"1900");
    gpmc_send('1',x"3009",x"0026");
    gpmc_send('1',x"300A",x"1A00");
    gpmc_send('1',x"300B",x"0025");
    gpmc_send('1',x"300C",x"1B00");
    gpmc_send('1',x"300D",x"0024");
    gpmc_send('1',x"300E",x"1C00");
    gpmc_send('1',x"300F",x"0023");
    gpmc_send('1',x"3010",x"1D00");
    gpmc_send('1',x"3011",x"0022");
    gpmc_send('1',x"3012",x"1E00");
    gpmc_send('1',x"3013",x"0021");
    gpmc_send('1',x"3014",x"1F00");
    gpmc_send('1',x"3015",x"0020");
    gpmc_send('1',x"3016",x"2000");
    gpmc_send('1',x"3017",x"001F");
    gpmc_send('1',x"3018",x"2100");
    gpmc_send('1',x"3019",x"001E");
    gpmc_send('1',x"301A",x"2200");
    gpmc_send('1',x"301B",x"001D");
    gpmc_send('1',x"301C",x"2300");
    gpmc_send('1',x"301D",x"001C");
    gpmc_send('1',x"301E",x"2400");
    gpmc_send('1',x"301F",x"001B");
    gpmc_send('1',x"3020",x"2500");
    gpmc_send('1',x"3021",x"001A");
    gpmc_send('1',x"3022",x"2600");
    gpmc_send('1',x"3023",x"0019");
    gpmc_send('1',x"3024",x"2700");
    gpmc_send('1',x"3025",x"0018");
    gpmc_send('1',x"3026",x"2800");
    gpmc_send('1',x"3027",x"0017");
    gpmc_send('1',x"3028",x"2900");
    gpmc_send('1',x"3029",x"0016");
    gpmc_send('1',x"302A",x"2A00");
    gpmc_send('1',x"302B",x"0015");
    gpmc_send('1',x"302C",x"2B00");
    gpmc_send('1',x"302D",x"0014");
    gpmc_send('1',x"302E",x"2C00");
    gpmc_send('1',x"302F",x"0013");
    gpmc_send('1',x"3030",x"2D00");
    gpmc_send('1',x"3031",x"0012");
    gpmc_send('1',x"3032",x"2E00");
    gpmc_send('1',x"3033",x"0011");
    gpmc_send('1',x"3034",x"2F00");
    gpmc_send('1',x"3035",x"0010");
    gpmc_send('1',x"3036",x"3000");
    gpmc_send('1',x"3037",x"000F");
    gpmc_send('1',x"3038",x"3100");
    gpmc_send('1',x"3039",x"000E");
    gpmc_send('1',x"303A",x"3200");
    gpmc_send('1',x"303B",x"000D");
    gpmc_send('1',x"303C",x"3300");
    gpmc_send('1',x"303D",x"000C");
    gpmc_send('1',x"303E",x"3400");
    gpmc_send('1',x"303F",x"000B");
    gpmc_send('1',x"3040",x"3500");
    gpmc_send('1',x"3041",x"000A");
    gpmc_send('1',x"3042",x"3600");
    gpmc_send('1',x"3043",x"0009");
    gpmc_send('1',x"3044",x"3700");
    gpmc_send('1',x"3045",x"0008");
    gpmc_send('1',x"3046",x"3800");
    gpmc_send('1',x"3047",x"0007");
    gpmc_send('1',x"3048",x"3900");
    gpmc_send('1',x"3049",x"0006");
    gpmc_send('1',x"304A",x"3A00");
    gpmc_send('1',x"304B",x"0005");
    gpmc_send('1',x"304C",x"3B00");
    gpmc_send('1',x"304D",x"0004");
    gpmc_send('1',x"304E",x"3C00");
    gpmc_send('1',x"304F",x"0003");
    gpmc_send('1',x"3050",x"3D00");
    gpmc_send('1',x"3051",x"0002");
    gpmc_send('1',x"3052",x"3E00");
    gpmc_send('1',x"3053",x"0001");
    gpmc_send('1',x"3054",x"3F00");
    gpmc_send('1',x"3055",x"0000");
    gpmc_send('1',x"3056",x"3F01");
    gpmc_send('1',x"3057",x"0000");
    gpmc_send('1',x"3058",x"3E02");
    gpmc_send('1',x"3059",x"0000");
    gpmc_send('1',x"305A",x"3D03");
    gpmc_send('1',x"305B",x"0000");
    gpmc_send('1',x"305C",x"3C04");
    gpmc_send('1',x"305D",x"0000");
    gpmc_send('1',x"305E",x"3B05");
    gpmc_send('1',x"305F",x"0000");
    gpmc_send('1',x"3060",x"3A06");
    gpmc_send('1',x"3061",x"0000");
    gpmc_send('1',x"3062",x"3907");
    gpmc_send('1',x"3063",x"0000");
    gpmc_send('1',x"3064",x"3808");
    gpmc_send('1',x"3065",x"0000");
    gpmc_send('1',x"3066",x"3709");
    gpmc_send('1',x"3067",x"0000");
    gpmc_send('1',x"3068",x"360A");
    gpmc_send('1',x"3069",x"0000");
    gpmc_send('1',x"306A",x"350B");
    gpmc_send('1',x"306B",x"0000");
    gpmc_send('1',x"306C",x"340C");
    gpmc_send('1',x"306D",x"0000");
    gpmc_send('1',x"306E",x"330D");
    gpmc_send('1',x"306F",x"0000");
    gpmc_send('1',x"3070",x"320E");
    gpmc_send('1',x"3071",x"0000");
    gpmc_send('1',x"3072",x"310F");
    gpmc_send('1',x"3073",x"0000");
    gpmc_send('1',x"3074",x"3010");
    gpmc_send('1',x"3075",x"0000");
    gpmc_send('1',x"3076",x"2F11");
    gpmc_send('1',x"3077",x"0000");
    gpmc_send('1',x"3078",x"2E12");
    gpmc_send('1',x"3079",x"0000");
    gpmc_send('1',x"307A",x"2D13");
    gpmc_send('1',x"307B",x"0000");
    gpmc_send('1',x"307C",x"2C14");
    gpmc_send('1',x"307D",x"0000");
    gpmc_send('1',x"307E",x"2B15");
    gpmc_send('1',x"307F",x"0000");
    gpmc_send('1',x"3080",x"2A16");
    gpmc_send('1',x"3081",x"0000");
    gpmc_send('1',x"3082",x"2917");
    gpmc_send('1',x"3083",x"0000");
    gpmc_send('1',x"3084",x"2818");
    gpmc_send('1',x"3085",x"0000");
    gpmc_send('1',x"3086",x"2719");
    gpmc_send('1',x"3087",x"0000");
    gpmc_send('1',x"3088",x"261A");
    gpmc_send('1',x"3089",x"0000");
    gpmc_send('1',x"308A",x"251B");
    gpmc_send('1',x"308B",x"0000");
    gpmc_send('1',x"308C",x"241C");
    gpmc_send('1',x"308D",x"0000");
    gpmc_send('1',x"308E",x"231D");
    gpmc_send('1',x"308F",x"0000");
    gpmc_send('1',x"3090",x"221E");
    gpmc_send('1',x"3091",x"0000");
    gpmc_send('1',x"3092",x"211F");
    gpmc_send('1',x"3093",x"0000");
    gpmc_send('1',x"3094",x"2020");
    gpmc_send('1',x"3095",x"0000");
    gpmc_send('1',x"3096",x"1F21");
    gpmc_send('1',x"3097",x"0000");
    gpmc_send('1',x"3098",x"1E22");
    gpmc_send('1',x"3099",x"0000");
    gpmc_send('1',x"309A",x"1D23");
    gpmc_send('1',x"309B",x"0000");
    gpmc_send('1',x"309C",x"1C24");
    gpmc_send('1',x"309D",x"0000");
    gpmc_send('1',x"309E",x"1B25");
    gpmc_send('1',x"309F",x"0000");
    gpmc_send('1',x"30A0",x"1A26");
    gpmc_send('1',x"30A1",x"0000");
    gpmc_send('1',x"30A2",x"1927");
    gpmc_send('1',x"30A3",x"0000");
    gpmc_send('1',x"30A4",x"1828");
    gpmc_send('1',x"30A5",x"0000");
    gpmc_send('1',x"30A6",x"1729");
    gpmc_send('1',x"30A7",x"0000");
    gpmc_send('1',x"30A8",x"162A");
    gpmc_send('1',x"30A9",x"0000");
    gpmc_send('1',x"30AA",x"152B");
    gpmc_send('1',x"30AB",x"0000");
    gpmc_send('1',x"30AC",x"142C");
    gpmc_send('1',x"30AD",x"0000");
    gpmc_send('1',x"30AE",x"132D");
    gpmc_send('1',x"30AF",x"0000");
    gpmc_send('1',x"30B0",x"122E");
    gpmc_send('1',x"30B1",x"0000");
    gpmc_send('1',x"30B2",x"112F");
    gpmc_send('1',x"30B3",x"0000");
    gpmc_send('1',x"30B4",x"1030");
    gpmc_send('1',x"30B5",x"0000");
    gpmc_send('1',x"30B6",x"0F31");
    gpmc_send('1',x"30B7",x"0000");
    gpmc_send('1',x"30B8",x"0E32");
    gpmc_send('1',x"30B9",x"0000");
    gpmc_send('1',x"30BA",x"0D33");
    gpmc_send('1',x"30BB",x"0000");
    gpmc_send('1',x"30BC",x"0C34");
    gpmc_send('1',x"30BD",x"0000");
    gpmc_send('1',x"30BE",x"0B35");
    gpmc_send('1',x"30BF",x"0000");
    gpmc_send('1',x"30C0",x"0A36");
    gpmc_send('1',x"30C1",x"0000");
    gpmc_send('1',x"30C2",x"0937");
    gpmc_send('1',x"30C3",x"0000");
    gpmc_send('1',x"30C4",x"0838");
    gpmc_send('1',x"30C5",x"0000");
    gpmc_send('1',x"30C6",x"0739");
    gpmc_send('1',x"30C7",x"0000");
    gpmc_send('1',x"30C8",x"063A");
    gpmc_send('1',x"30C9",x"0000");
    gpmc_send('1',x"30CA",x"053B");
    gpmc_send('1',x"30CB",x"0000");
    gpmc_send('1',x"30CC",x"043C");
    gpmc_send('1',x"30CD",x"0000");
    gpmc_send('1',x"30CE",x"033D");
    gpmc_send('1',x"30CF",x"0000");
    gpmc_send('1',x"30D0",x"023E");
    gpmc_send('1',x"30D1",x"0000");
    gpmc_send('1',x"30D2",x"013F");
    gpmc_send('1',x"30D3",x"0000");
    gpmc_send('1',x"30D4",x"003F");
    gpmc_send('1',x"30D5",x"0000");
    gpmc_send('1',x"30D6",x"003E");
    gpmc_send('1',x"30D7",x"0001");
    gpmc_send('1',x"30D8",x"003D");
    gpmc_send('1',x"30D9",x"0002");
    gpmc_send('1',x"30DA",x"003C");
    gpmc_send('1',x"30DB",x"0003");
    gpmc_send('1',x"30DC",x"003B");
    gpmc_send('1',x"30DD",x"0004");
    gpmc_send('1',x"30DE",x"003A");
    gpmc_send('1',x"30DF",x"0005");
    gpmc_send('1',x"30E0",x"0039");
    gpmc_send('1',x"30E1",x"0006");
    gpmc_send('1',x"30E2",x"0038");
    gpmc_send('1',x"30E3",x"0007");
    gpmc_send('1',x"30E4",x"0037");
    gpmc_send('1',x"30E5",x"0008");
    gpmc_send('1',x"30E6",x"0036");
    gpmc_send('1',x"30E7",x"0009");
    gpmc_send('1',x"30E8",x"0035");
    gpmc_send('1',x"30E9",x"000A");
    gpmc_send('1',x"30EA",x"0034");
    gpmc_send('1',x"30EB",x"000B");
    gpmc_send('1',x"30EC",x"0033");
    gpmc_send('1',x"30ED",x"000C");
    gpmc_send('1',x"30EE",x"0032");
    gpmc_send('1',x"30EF",x"000D");
    gpmc_send('1',x"30F0",x"0031");
    gpmc_send('1',x"30F1",x"000E");
    gpmc_send('1',x"30F2",x"0030");
    gpmc_send('1',x"30F3",x"000F");
    gpmc_send('1',x"30F4",x"002F");
    gpmc_send('1',x"30F5",x"0010");
    gpmc_send('1',x"30F6",x"002E");
    gpmc_send('1',x"30F7",x"0011");
    gpmc_send('1',x"30F8",x"002D");
    gpmc_send('1',x"30F9",x"0012");
    gpmc_send('1',x"30FA",x"002C");
    gpmc_send('1',x"30FB",x"0013");
    gpmc_send('1',x"30FC",x"002B");
    gpmc_send('1',x"30FD",x"0014");
    gpmc_send('1',x"30FE",x"002A");
    gpmc_send('1',x"30FF",x"0015");
    gpmc_send('1',x"3100",x"0029");
    gpmc_send('1',x"3101",x"0016");
    gpmc_send('1',x"3102",x"0028");
    gpmc_send('1',x"3103",x"0017");
    gpmc_send('1',x"3104",x"0027");
    gpmc_send('1',x"3105",x"0018");
    gpmc_send('1',x"3106",x"0026");
    gpmc_send('1',x"3107",x"0019");
    gpmc_send('1',x"3108",x"0025");
    gpmc_send('1',x"3109",x"001A");
    gpmc_send('1',x"310A",x"0024");
    gpmc_send('1',x"310B",x"001B");
    gpmc_send('1',x"310C",x"0023");
    gpmc_send('1',x"310D",x"001C");
    gpmc_send('1',x"310E",x"0022");
    gpmc_send('1',x"310F",x"001D");
    gpmc_send('1',x"3110",x"0021");
    gpmc_send('1',x"3111",x"001E");
    gpmc_send('1',x"3112",x"0020");
    gpmc_send('1',x"3113",x"001F");
    gpmc_send('1',x"3114",x"001F");
    gpmc_send('1',x"3115",x"0020");
    gpmc_send('1',x"3116",x"001E");
    gpmc_send('1',x"3117",x"0021");
    gpmc_send('1',x"3118",x"001D");
    gpmc_send('1',x"3119",x"0022");
    gpmc_send('1',x"311A",x"001C");
    gpmc_send('1',x"311B",x"0023");
    gpmc_send('1',x"311C",x"001B");
    gpmc_send('1',x"311D",x"0024");
    gpmc_send('1',x"311E",x"001A");
    gpmc_send('1',x"311F",x"0025");
    gpmc_send('1',x"3120",x"0019");
    gpmc_send('1',x"3121",x"0026");
    gpmc_send('1',x"3122",x"0018");
    gpmc_send('1',x"3123",x"0027");
    gpmc_send('1',x"3124",x"0017");
    gpmc_send('1',x"3125",x"0028");
    gpmc_send('1',x"3126",x"0016");
    gpmc_send('1',x"3127",x"0029");
    gpmc_send('1',x"3128",x"0015");
    gpmc_send('1',x"3129",x"002A");
    gpmc_send('1',x"312A",x"0014");
    gpmc_send('1',x"312B",x"002B");
    gpmc_send('1',x"312C",x"0013");
    gpmc_send('1',x"312D",x"002C");
    gpmc_send('1',x"312E",x"0012");
    gpmc_send('1',x"312F",x"002D");
    gpmc_send('1',x"3130",x"0011");
    gpmc_send('1',x"3131",x"002E");
    gpmc_send('1',x"3132",x"0010");
    gpmc_send('1',x"3133",x"002F");
    gpmc_send('1',x"3134",x"000F");
    gpmc_send('1',x"3135",x"0030");
    gpmc_send('1',x"3136",x"000E");
    gpmc_send('1',x"3137",x"0031");
    gpmc_send('1',x"3138",x"000D");
    gpmc_send('1',x"3139",x"0032");
    gpmc_send('1',x"313A",x"000C");
    gpmc_send('1',x"313B",x"0033");
    gpmc_send('1',x"313C",x"000B");
    gpmc_send('1',x"313D",x"0034");
    gpmc_send('1',x"313E",x"000A");
    gpmc_send('1',x"313F",x"0035");
    gpmc_send('1',x"3140",x"0009");
    gpmc_send('1',x"3141",x"0036");
    gpmc_send('1',x"3142",x"0008");
    gpmc_send('1',x"3143",x"0037");
    gpmc_send('1',x"3144",x"0007");
    gpmc_send('1',x"3145",x"0038");
    gpmc_send('1',x"3146",x"0006");
    gpmc_send('1',x"3147",x"0039");
    gpmc_send('1',x"3148",x"0005");
    gpmc_send('1',x"3149",x"003A");
    gpmc_send('1',x"314A",x"0004");
    gpmc_send('1',x"314B",x"003B");
    gpmc_send('1',x"314C",x"0003");
    gpmc_send('1',x"314D",x"003C");
    gpmc_send('1',x"314E",x"0002");
    gpmc_send('1',x"314F",x"003D");
    gpmc_send('1',x"3150",x"0001");
    gpmc_send('1',x"3151",x"003E");
    gpmc_send('1',x"3152",x"0000");
    gpmc_send('1',x"3153",x"003F");
    gpmc_send('1',x"3154",x"0100");
    gpmc_send('1',x"3155",x"003E");
    gpmc_send('1',x"3156",x"0200");
    gpmc_send('1',x"3157",x"003D");
    gpmc_send('1',x"3158",x"0300");
    gpmc_send('1',x"3159",x"003C");
    gpmc_send('1',x"315A",x"0400");
    gpmc_send('1',x"315B",x"003B");
    gpmc_send('1',x"315C",x"0500");
    gpmc_send('1',x"315D",x"003A");
    gpmc_send('1',x"315E",x"0600");
    gpmc_send('1',x"315F",x"0039");
    gpmc_send('1',x"3160",x"0700");
    gpmc_send('1',x"3161",x"0038");
    gpmc_send('1',x"3162",x"0800");
    gpmc_send('1',x"3163",x"0037");
    gpmc_send('1',x"3164",x"0900");
    gpmc_send('1',x"3165",x"0036");
    gpmc_send('1',x"3166",x"0A00");
    gpmc_send('1',x"3167",x"0035");
    gpmc_send('1',x"3168",x"0B00");
    gpmc_send('1',x"3169",x"0034");
    gpmc_send('1',x"316A",x"0C00");
    gpmc_send('1',x"316B",x"0033");
    gpmc_send('1',x"316C",x"0D00");
    gpmc_send('1',x"316D",x"0032");
    gpmc_send('1',x"316E",x"0E00");
    gpmc_send('1',x"316F",x"0031");
    gpmc_send('1',x"3170",x"0F00");
    gpmc_send('1',x"3171",x"0030");
    gpmc_send('1',x"3172",x"1000");
    gpmc_send('1',x"3173",x"002F");
    gpmc_send('1',x"3174",x"1100");
    gpmc_send('1',x"3175",x"002E");
    gpmc_send('1',x"3176",x"1200");
    gpmc_send('1',x"3177",x"002D");
    gpmc_send('1',x"3178",x"1300");
    gpmc_send('1',x"3179",x"002C");
    gpmc_send('1',x"317A",x"1400");
    gpmc_send('1',x"317B",x"002B");
    gpmc_send('1',x"317C",x"1500");
    gpmc_send('1',x"317D",x"002A");
    gpmc_send('1',x"317E",x"1600");
    gpmc_send('1',x"317F",x"0029");
    gpmc_send('1',x"3180",x"1700");
    gpmc_send('1',x"3181",x"0028");
    gpmc_send('1',x"3182",x"1800");
    gpmc_send('1',x"3183",x"0027");
    gpmc_send('1',x"3184",x"1900");
    gpmc_send('1',x"3185",x"0026");
    gpmc_send('1',x"3186",x"1A00");
    gpmc_send('1',x"3187",x"0025");
    gpmc_send('1',x"3188",x"1B00");
    gpmc_send('1',x"3189",x"0024");
    gpmc_send('1',x"318A",x"1C00");
    gpmc_send('1',x"318B",x"0023");
    gpmc_send('1',x"318C",x"1D00");
    gpmc_send('1',x"318D",x"0022");
    gpmc_send('1',x"318E",x"1E00");
    gpmc_send('1',x"318F",x"0021");
    gpmc_send('1',x"3190",x"1F00");
    gpmc_send('1',x"3191",x"0020");
    gpmc_send('1',x"3192",x"2000");
    gpmc_send('1',x"3193",x"001F");
    gpmc_send('1',x"3194",x"2100");
    gpmc_send('1',x"3195",x"001E");
    gpmc_send('1',x"3196",x"2200");
    gpmc_send('1',x"3197",x"001D");
    gpmc_send('1',x"3198",x"2300");
    gpmc_send('1',x"3199",x"001C");
    gpmc_send('1',x"319A",x"2400");
    gpmc_send('1',x"319B",x"001B");
    gpmc_send('1',x"319C",x"2500");
    gpmc_send('1',x"319D",x"001A");
    gpmc_send('1',x"319E",x"2600");
    gpmc_send('1',x"319F",x"0019");
    gpmc_send('1',x"31A0",x"2700");
    gpmc_send('1',x"31A1",x"0018");
    gpmc_send('1',x"31A2",x"2800");
    gpmc_send('1',x"31A3",x"0017");
    gpmc_send('1',x"31A4",x"2900");
    gpmc_send('1',x"31A5",x"0016");
    gpmc_send('1',x"31A6",x"2A00");
    gpmc_send('1',x"31A7",x"0015");
    gpmc_send('1',x"31A8",x"2B00");
    gpmc_send('1',x"31A9",x"0014");
    gpmc_send('1',x"31AA",x"2C00");
    gpmc_send('1',x"31AB",x"0013");
    gpmc_send('1',x"31AC",x"2D00");
    gpmc_send('1',x"31AD",x"0012");
    gpmc_send('1',x"31AE",x"2E00");
    gpmc_send('1',x"31AF",x"0011");
    gpmc_send('1',x"31B0",x"2F00");
    gpmc_send('1',x"31B1",x"0010");
    gpmc_send('1',x"31B2",x"3000");
    gpmc_send('1',x"31B3",x"000F");
    gpmc_send('1',x"31B4",x"3100");
    gpmc_send('1',x"31B5",x"000E");
    gpmc_send('1',x"31B6",x"3200");
    gpmc_send('1',x"31B7",x"000D");
    gpmc_send('1',x"31B8",x"3300");
    gpmc_send('1',x"31B9",x"000C");
    gpmc_send('1',x"31BA",x"3400");
    gpmc_send('1',x"31BB",x"000B");
    gpmc_send('1',x"31BC",x"3500");
    gpmc_send('1',x"31BD",x"000A");
    gpmc_send('1',x"31BE",x"3600");
    gpmc_send('1',x"31BF",x"0009");
    gpmc_send('1',x"31C0",x"3700");
    gpmc_send('1',x"31C1",x"0008");
    gpmc_send('1',x"31C2",x"3800");
    gpmc_send('1',x"31C3",x"0007");
    gpmc_send('1',x"31C4",x"3900");
    gpmc_send('1',x"31C5",x"0006");
    gpmc_send('1',x"31C6",x"3A00");
    gpmc_send('1',x"31C7",x"0005");
    gpmc_send('1',x"31C8",x"3B00");
    gpmc_send('1',x"31C9",x"0004");
    gpmc_send('1',x"31CA",x"3C00");
    gpmc_send('1',x"31CB",x"0003");
    gpmc_send('1',x"31CC",x"3D00");
    gpmc_send('1',x"31CD",x"0002");
    gpmc_send('1',x"31CE",x"3E00");
    gpmc_send('1',x"31CF",x"0001");
    gpmc_send('1',x"31D0",x"3F00");
    gpmc_send('1',x"31D1",x"0000");
    gpmc_send('1',x"31D2",x"3F01");
    gpmc_send('1',x"31D3",x"0000");
    gpmc_send('1',x"31D4",x"3E02");
    gpmc_send('1',x"31D5",x"0000");
    gpmc_send('1',x"31D6",x"3D03");
    gpmc_send('1',x"31D7",x"0000");
    gpmc_send('1',x"31D8",x"3C04");
    gpmc_send('1',x"31D9",x"0000");
    gpmc_send('1',x"31DA",x"3B05");
    gpmc_send('1',x"31DB",x"0000");
    gpmc_send('1',x"31DC",x"3A06");
    gpmc_send('1',x"31DD",x"0000");
    gpmc_send('1',x"31DE",x"3907");
    gpmc_send('1',x"31DF",x"0000");
    gpmc_send('1',x"31E0",x"3808");
    gpmc_send('1',x"31E1",x"0000");
    gpmc_send('1',x"31E2",x"3709");
    gpmc_send('1',x"31E3",x"0000");
    gpmc_send('1',x"31E4",x"360A");
    gpmc_send('1',x"31E5",x"0000");
    gpmc_send('1',x"31E6",x"350B");
    gpmc_send('1',x"31E7",x"0000");
    gpmc_send('1',x"31E8",x"340C");
    gpmc_send('1',x"31E9",x"0000");
    gpmc_send('1',x"31EA",x"330D");
    gpmc_send('1',x"31EB",x"0000");
    gpmc_send('1',x"31EC",x"320E");
    gpmc_send('1',x"31ED",x"0000");
    gpmc_send('1',x"31EE",x"310F");
    gpmc_send('1',x"31EF",x"0000");
    gpmc_send('1',x"31F0",x"3010");
    gpmc_send('1',x"31F1",x"0000");
    gpmc_send('1',x"31F2",x"2F11");
    gpmc_send('1',x"31F3",x"0000");
    gpmc_send('1',x"31F4",x"2E12");
    gpmc_send('1',x"31F5",x"0000");
    gpmc_send('1',x"31F6",x"2D13");
    gpmc_send('1',x"31F7",x"0000");
    gpmc_send('1',x"31F8",x"2C14");
    gpmc_send('1',x"31F9",x"0000");
    gpmc_send('1',x"31FA",x"2B15");
    gpmc_send('1',x"31FB",x"0000");
    gpmc_send('1',x"31FC",x"2A16");
    gpmc_send('1',x"31FD",x"0000");
    gpmc_send('1',x"31FE",x"2917");
    gpmc_send('1',x"31FF",x"0000");
    gpmc_send('1',x"3200",x"2818");
    gpmc_send('1',x"3201",x"0000");
    gpmc_send('1',x"3202",x"2719");
    gpmc_send('1',x"3203",x"0000");
    gpmc_send('1',x"3204",x"261A");
    gpmc_send('1',x"3205",x"0000");
    gpmc_send('1',x"3206",x"251B");
    gpmc_send('1',x"3207",x"0000");
    gpmc_send('1',x"3208",x"241C");
    gpmc_send('1',x"3209",x"0000");
    gpmc_send('1',x"320A",x"231D");
    gpmc_send('1',x"320B",x"0000");
    gpmc_send('1',x"320C",x"221E");
    gpmc_send('1',x"320D",x"0000");
    gpmc_send('1',x"320E",x"211F");
    gpmc_send('1',x"320F",x"0000");
    gpmc_send('1',x"3210",x"2020");
    gpmc_send('1',x"3211",x"0000");
    gpmc_send('1',x"3212",x"1F21");
    gpmc_send('1',x"3213",x"0000");
    gpmc_send('1',x"3214",x"1E22");
    gpmc_send('1',x"3215",x"0000");
    gpmc_send('1',x"3216",x"1D23");
    gpmc_send('1',x"3217",x"0000");
    gpmc_send('1',x"3218",x"1C24");
    gpmc_send('1',x"3219",x"0000");
    gpmc_send('1',x"321A",x"1B25");
    gpmc_send('1',x"321B",x"0000");
    gpmc_send('1',x"321C",x"1A26");
    gpmc_send('1',x"321D",x"0000");
    gpmc_send('1',x"321E",x"1927");
    gpmc_send('1',x"321F",x"0000");
    gpmc_send('1',x"3220",x"1828");
    gpmc_send('1',x"3221",x"0000");
    gpmc_send('1',x"3222",x"1729");
    gpmc_send('1',x"3223",x"0000");
    gpmc_send('1',x"3224",x"162A");
    gpmc_send('1',x"3225",x"0000");
    gpmc_send('1',x"3226",x"152B");
    gpmc_send('1',x"3227",x"0000");
    gpmc_send('1',x"3228",x"142C");
    gpmc_send('1',x"3229",x"0000");
    gpmc_send('1',x"322A",x"132D");
    gpmc_send('1',x"322B",x"0000");
    gpmc_send('1',x"322C",x"122E");
    gpmc_send('1',x"322D",x"0000");
    gpmc_send('1',x"322E",x"112F");
    gpmc_send('1',x"322F",x"0000");
    gpmc_send('1',x"3230",x"1030");
    gpmc_send('1',x"3231",x"0000");
    gpmc_send('1',x"3232",x"0F31");
    gpmc_send('1',x"3233",x"0000");
    gpmc_send('1',x"3234",x"0E32");
    gpmc_send('1',x"3235",x"0000");
    gpmc_send('1',x"3236",x"0D33");
    gpmc_send('1',x"3237",x"0000");
    gpmc_send('1',x"3238",x"0C34");
    gpmc_send('1',x"3239",x"0000");
    gpmc_send('1',x"323A",x"0B35");
    gpmc_send('1',x"323B",x"0000");
    gpmc_send('1',x"323C",x"0A36");
    gpmc_send('1',x"323D",x"0000");
    gpmc_send('1',x"323E",x"0937");
    gpmc_send('1',x"323F",x"0000");
    gpmc_send('1',x"3240",x"0838");
    gpmc_send('1',x"3241",x"0000");
    gpmc_send('1',x"3242",x"0739");
    gpmc_send('1',x"3243",x"0000");
    gpmc_send('1',x"3244",x"063A");
    gpmc_send('1',x"3245",x"0000");
    gpmc_send('1',x"3246",x"053B");
    gpmc_send('1',x"3247",x"0000");
    gpmc_send('1',x"3248",x"043C");
    gpmc_send('1',x"3249",x"0000");
    gpmc_send('1',x"324A",x"033D");
    gpmc_send('1',x"324B",x"0000");
    gpmc_send('1',x"324C",x"023E");
    gpmc_send('1',x"324D",x"0000");
    gpmc_send('1',x"324E",x"013F");
    gpmc_send('1',x"324F",x"0000");
    gpmc_send('1',x"3250",x"003F");
    gpmc_send('1',x"3251",x"0000");
    gpmc_send('1',x"3252",x"003E");
    gpmc_send('1',x"3253",x"0001");
    gpmc_send('1',x"3254",x"003D");
    gpmc_send('1',x"3255",x"0002");
    gpmc_send('1',x"3256",x"003C");
    gpmc_send('1',x"3257",x"0003");
    gpmc_send('1',x"3258",x"003B");
    gpmc_send('1',x"3259",x"0004");
    gpmc_send('1',x"325A",x"003A");
    gpmc_send('1',x"325B",x"0005");
    gpmc_send('1',x"325C",x"0039");
    gpmc_send('1',x"325D",x"0006");
    gpmc_send('1',x"325E",x"0038");
    gpmc_send('1',x"325F",x"0007");
    gpmc_send('1',x"3260",x"0037");
    gpmc_send('1',x"3261",x"0008");
    gpmc_send('1',x"3262",x"0036");
    gpmc_send('1',x"3263",x"0009");
    gpmc_send('1',x"3264",x"0035");
    gpmc_send('1',x"3265",x"000A");
    gpmc_send('1',x"3266",x"0034");
    gpmc_send('1',x"3267",x"000B");
    gpmc_send('1',x"3268",x"0033");
    gpmc_send('1',x"3269",x"000C");
    gpmc_send('1',x"326A",x"0032");
    gpmc_send('1',x"326B",x"000D");
    gpmc_send('1',x"326C",x"0031");
    gpmc_send('1',x"326D",x"000E");
    gpmc_send('1',x"326E",x"0030");
    gpmc_send('1',x"326F",x"000F");
    gpmc_send('1',x"3270",x"002F");
    gpmc_send('1',x"3271",x"0010");
    gpmc_send('1',x"3272",x"002E");
    gpmc_send('1',x"3273",x"0011");
    gpmc_send('1',x"3274",x"002D");
    gpmc_send('1',x"3275",x"0012");
    gpmc_send('1',x"3276",x"002C");
    gpmc_send('1',x"3277",x"0013");
    gpmc_send('1',x"3278",x"002B");
    gpmc_send('1',x"3279",x"0014");
    gpmc_send('1',x"327A",x"002A");
    gpmc_send('1',x"327B",x"0015");
    gpmc_send('1',x"327C",x"0029");
    gpmc_send('1',x"327D",x"0016");
    gpmc_send('1',x"327E",x"0028");
    gpmc_send('1',x"327F",x"0017");
    gpmc_send('1',x"3280",x"0027");
    gpmc_send('1',x"3281",x"0018");
    gpmc_send('1',x"3282",x"0026");
    gpmc_send('1',x"3283",x"0019");
    gpmc_send('1',x"3284",x"0025");
    gpmc_send('1',x"3285",x"001A");
    gpmc_send('1',x"3286",x"0024");
    gpmc_send('1',x"3287",x"001B");
    gpmc_send('1',x"3288",x"0023");
    gpmc_send('1',x"3289",x"001C");
    gpmc_send('1',x"328A",x"0022");
    gpmc_send('1',x"328B",x"001D");
    gpmc_send('1',x"328C",x"0021");
    gpmc_send('1',x"328D",x"001E");
    gpmc_send('1',x"328E",x"0020");
    gpmc_send('1',x"328F",x"001F");
    gpmc_send('1',x"3290",x"001F");
    gpmc_send('1',x"3291",x"0020");
    gpmc_send('1',x"3292",x"001E");
    gpmc_send('1',x"3293",x"0021");
    gpmc_send('1',x"3294",x"001D");
    gpmc_send('1',x"3295",x"0022");
    gpmc_send('1',x"3296",x"001C");
    gpmc_send('1',x"3297",x"0023");
    gpmc_send('1',x"3298",x"001B");
    gpmc_send('1',x"3299",x"0024");
    gpmc_send('1',x"329A",x"001A");
    gpmc_send('1',x"329B",x"0025");
    gpmc_send('1',x"329C",x"0019");
    gpmc_send('1',x"329D",x"0026");
    gpmc_send('1',x"329E",x"0018");
    gpmc_send('1',x"329F",x"0027");
    gpmc_send('1',x"32A0",x"0017");
    gpmc_send('1',x"32A1",x"0028");
    gpmc_send('1',x"32A2",x"0016");
    gpmc_send('1',x"32A3",x"0029");
    gpmc_send('1',x"32A4",x"0015");
    gpmc_send('1',x"32A5",x"002A");
    gpmc_send('1',x"32A6",x"0014");
    gpmc_send('1',x"32A7",x"002B");
    gpmc_send('1',x"32A8",x"0013");
    gpmc_send('1',x"32A9",x"002C");
    gpmc_send('1',x"32AA",x"0012");
    gpmc_send('1',x"32AB",x"002D");
    gpmc_send('1',x"32AC",x"0011");
    gpmc_send('1',x"32AD",x"002E");
    gpmc_send('1',x"32AE",x"0010");
    gpmc_send('1',x"32AF",x"002F");
    gpmc_send('1',x"32B0",x"000F");
    gpmc_send('1',x"32B1",x"0030");
    gpmc_send('1',x"32B2",x"000E");
    gpmc_send('1',x"32B3",x"0031");
    gpmc_send('1',x"32B4",x"000D");
    gpmc_send('1',x"32B5",x"0032");
    gpmc_send('1',x"32B6",x"000C");
    gpmc_send('1',x"32B7",x"0033");
    gpmc_send('1',x"32B8",x"000B");
    gpmc_send('1',x"32B9",x"0034");
    gpmc_send('1',x"32BA",x"000A");
    gpmc_send('1',x"32BB",x"0035");
    gpmc_send('1',x"32BC",x"0009");
    gpmc_send('1',x"32BD",x"0036");
    gpmc_send('1',x"32BE",x"0008");
    gpmc_send('1',x"32BF",x"0037");
    gpmc_send('1',x"32C0",x"0007");
    gpmc_send('1',x"32C1",x"0038");
    gpmc_send('1',x"32C2",x"0006");
    gpmc_send('1',x"32C3",x"0039");
    gpmc_send('1',x"32C4",x"0005");
    gpmc_send('1',x"32C5",x"003A");
    gpmc_send('1',x"32C6",x"0004");
    gpmc_send('1',x"32C7",x"003B");
    gpmc_send('1',x"32C8",x"0003");
    gpmc_send('1',x"32C9",x"003C");
    gpmc_send('1',x"32CA",x"0002");
    gpmc_send('1',x"32CB",x"003D");
    gpmc_send('1',x"32CC",x"0001");
    gpmc_send('1',x"32CD",x"003E");
    gpmc_send('1',x"32CE",x"0000");
    gpmc_send('1',x"32CF",x"003F");
    gpmc_send('1',x"32D0",x"0100");
    gpmc_send('1',x"32D1",x"003E");
    gpmc_send('1',x"32D2",x"0200");
    gpmc_send('1',x"32D3",x"003D");
    gpmc_send('1',x"32D4",x"0300");
    gpmc_send('1',x"32D5",x"003C");
    gpmc_send('1',x"32D6",x"0400");
    gpmc_send('1',x"32D7",x"003B");
    gpmc_send('1',x"32D8",x"0500");
    gpmc_send('1',x"32D9",x"003A");
    gpmc_send('1',x"32DA",x"0600");
    gpmc_send('1',x"32DB",x"0039");
    gpmc_send('1',x"32DC",x"0700");
    gpmc_send('1',x"32DD",x"0038");
    gpmc_send('1',x"32DE",x"0800");
    gpmc_send('1',x"32DF",x"0037");
    gpmc_send('1',x"32E0",x"0900");
    gpmc_send('1',x"32E1",x"0036");
    gpmc_send('1',x"32E2",x"0A00");
    gpmc_send('1',x"32E3",x"0035");
    gpmc_send('1',x"32E4",x"0B00");
    gpmc_send('1',x"32E5",x"0034");
    gpmc_send('1',x"32E6",x"0C00");
    gpmc_send('1',x"32E7",x"0033");
    gpmc_send('1',x"32E8",x"0D00");
    gpmc_send('1',x"32E9",x"0032");
    gpmc_send('1',x"32EA",x"0E00");
    gpmc_send('1',x"32EB",x"0031");
    gpmc_send('1',x"32EC",x"0F00");
    gpmc_send('1',x"32ED",x"0030");
    gpmc_send('1',x"32EE",x"1000");
    gpmc_send('1',x"32EF",x"002F");
    gpmc_send('1',x"32F0",x"1100");
    gpmc_send('1',x"32F1",x"002E");
    gpmc_send('1',x"32F2",x"1200");
    gpmc_send('1',x"32F3",x"002D");
    gpmc_send('1',x"32F4",x"1300");
    gpmc_send('1',x"32F5",x"002C");
    gpmc_send('1',x"32F6",x"1400");
    gpmc_send('1',x"32F7",x"002B");
    gpmc_send('1',x"32F8",x"1500");
    gpmc_send('1',x"32F9",x"002A");
    gpmc_send('1',x"32FA",x"1600");
    gpmc_send('1',x"32FB",x"0029");
    gpmc_send('1',x"32FC",x"1700");
    gpmc_send('1',x"32FD",x"0028");
    gpmc_send('1',x"32FE",x"1800");
    gpmc_send('1',x"32FF",x"0027");
    gpmc_send('1',x"3300",x"1900");
    gpmc_send('1',x"3301",x"0026");
    gpmc_send('1',x"3302",x"1A00");
    gpmc_send('1',x"3303",x"0025");
    gpmc_send('1',x"3304",x"1B00");
    gpmc_send('1',x"3305",x"0024");
    gpmc_send('1',x"3306",x"1C00");
    gpmc_send('1',x"3307",x"0023");
    gpmc_send('1',x"3308",x"1D00");
    gpmc_send('1',x"3309",x"0022");
    gpmc_send('1',x"330A",x"1E00");
    gpmc_send('1',x"330B",x"0021");
    gpmc_send('1',x"330C",x"1F00");
    gpmc_send('1',x"330D",x"0020");
    gpmc_send('1',x"330E",x"2000");
    gpmc_send('1',x"330F",x"001F");
    gpmc_send('1',x"3310",x"2100");
    gpmc_send('1',x"3311",x"001E");
    gpmc_send('1',x"3312",x"2200");
    gpmc_send('1',x"3313",x"001D");
    gpmc_send('1',x"3314",x"2300");
    gpmc_send('1',x"3315",x"001C");
    gpmc_send('1',x"3316",x"2400");
    gpmc_send('1',x"3317",x"001B");
    gpmc_send('1',x"3318",x"2500");
    gpmc_send('1',x"3319",x"001A");
    gpmc_send('1',x"331A",x"2600");
    gpmc_send('1',x"331B",x"0019");
    gpmc_send('1',x"331C",x"2700");
    gpmc_send('1',x"331D",x"0018");
    gpmc_send('1',x"331E",x"2800");
    gpmc_send('1',x"331F",x"0017");
    gpmc_send('1',x"3320",x"2900");
    gpmc_send('1',x"3321",x"0016");
    gpmc_send('1',x"3322",x"2A00");
    gpmc_send('1',x"3323",x"0015");
    gpmc_send('1',x"3324",x"2B00");
    gpmc_send('1',x"3325",x"0014");
    gpmc_send('1',x"3326",x"2C00");
    gpmc_send('1',x"3327",x"0013");
    gpmc_send('1',x"3328",x"2D00");
    gpmc_send('1',x"3329",x"0012");
    gpmc_send('1',x"332A",x"2E00");
    gpmc_send('1',x"332B",x"0011");
    gpmc_send('1',x"332C",x"2F00");
    gpmc_send('1',x"332D",x"0010");
    gpmc_send('1',x"332E",x"3000");
    gpmc_send('1',x"332F",x"000F");
    gpmc_send('1',x"3330",x"3100");
    gpmc_send('1',x"3331",x"000E");
    gpmc_send('1',x"3332",x"3200");
    gpmc_send('1',x"3333",x"000D");
    gpmc_send('1',x"3334",x"3300");
    gpmc_send('1',x"3335",x"000C");
    gpmc_send('1',x"3336",x"3400");
    gpmc_send('1',x"3337",x"000B");
    gpmc_send('1',x"3338",x"3500");
    gpmc_send('1',x"3339",x"000A");
    gpmc_send('1',x"333A",x"3600");
    gpmc_send('1',x"333B",x"0009");
    gpmc_send('1',x"333C",x"3700");
    gpmc_send('1',x"333D",x"0008");
    gpmc_send('1',x"333E",x"3800");
    gpmc_send('1',x"333F",x"0007");
    gpmc_send('1',x"3340",x"3900");
    gpmc_send('1',x"3341",x"0006");
    gpmc_send('1',x"3342",x"3A00");
    gpmc_send('1',x"3343",x"0005");
    gpmc_send('1',x"3344",x"3B00");
    gpmc_send('1',x"3345",x"0004");
    gpmc_send('1',x"3346",x"3C00");
    gpmc_send('1',x"3347",x"0003");
    gpmc_send('1',x"3348",x"3D00");
    gpmc_send('1',x"3349",x"0002");
    gpmc_send('1',x"334A",x"3E00");
    gpmc_send('1',x"334B",x"0001");
    gpmc_send('1',x"334C",x"3F00");
    gpmc_send('1',x"334D",x"0000");
    gpmc_send('1',x"334E",x"3F01");
    gpmc_send('1',x"334F",x"0000");
    gpmc_send('1',x"3350",x"3E02");
    gpmc_send('1',x"3351",x"0000");
    gpmc_send('1',x"3352",x"3D03");
    gpmc_send('1',x"3353",x"0000");
    gpmc_send('1',x"3354",x"3C04");
    gpmc_send('1',x"3355",x"0000");
    gpmc_send('1',x"3356",x"3B05");
    gpmc_send('1',x"3357",x"0000");
    gpmc_send('1',x"3358",x"3A06");
    gpmc_send('1',x"3359",x"0000");
    gpmc_send('1',x"335A",x"3907");
    gpmc_send('1',x"335B",x"0000");
    gpmc_send('1',x"335C",x"3808");
    gpmc_send('1',x"335D",x"0000");
    gpmc_send('1',x"335E",x"3709");
    gpmc_send('1',x"335F",x"0000");
    gpmc_send('1',x"3360",x"360A");
    gpmc_send('1',x"3361",x"0000");
    gpmc_send('1',x"3362",x"350B");
    gpmc_send('1',x"3363",x"0000");
    gpmc_send('1',x"3364",x"340C");
    gpmc_send('1',x"3365",x"0000");
    gpmc_send('1',x"3366",x"330D");
    gpmc_send('1',x"3367",x"0000");
    gpmc_send('1',x"3368",x"320E");
    gpmc_send('1',x"3369",x"0000");
    gpmc_send('1',x"336A",x"310F");
    gpmc_send('1',x"336B",x"0000");
    gpmc_send('1',x"336C",x"3010");
    gpmc_send('1',x"336D",x"0000");
    gpmc_send('1',x"336E",x"2F11");
    gpmc_send('1',x"336F",x"0000");
    gpmc_send('1',x"3370",x"2E12");
    gpmc_send('1',x"3371",x"0000");
    gpmc_send('1',x"3372",x"2D13");
    gpmc_send('1',x"3373",x"0000");
    gpmc_send('1',x"3374",x"2C14");
    gpmc_send('1',x"3375",x"0000");
    gpmc_send('1',x"3376",x"2B15");
    gpmc_send('1',x"3377",x"0000");
    gpmc_send('1',x"3378",x"2A16");
    gpmc_send('1',x"3379",x"0000");
    gpmc_send('1',x"337A",x"2917");
    gpmc_send('1',x"337B",x"0000");
    gpmc_send('1',x"337C",x"2818");
    gpmc_send('1',x"337D",x"0000");
    gpmc_send('1',x"337E",x"2719");
    gpmc_send('1',x"337F",x"0000");
    gpmc_send('1',x"3380",x"261A");
    gpmc_send('1',x"3381",x"0000");
    gpmc_send('1',x"3382",x"251B");
    gpmc_send('1',x"3383",x"0000");
    gpmc_send('1',x"3384",x"241C");
    gpmc_send('1',x"3385",x"0000");
    gpmc_send('1',x"3386",x"231D");
    gpmc_send('1',x"3387",x"0000");
    gpmc_send('1',x"3388",x"221E");
    gpmc_send('1',x"3389",x"0000");
    gpmc_send('1',x"338A",x"211F");
    gpmc_send('1',x"338B",x"0000");
    gpmc_send('1',x"338C",x"2020");
    gpmc_send('1',x"338D",x"0000");
    gpmc_send('1',x"338E",x"1F21");
    gpmc_send('1',x"338F",x"0000");
    gpmc_send('1',x"3390",x"1E22");
    gpmc_send('1',x"3391",x"0000");
    gpmc_send('1',x"3392",x"1D23");
    gpmc_send('1',x"3393",x"0000");
    gpmc_send('1',x"3394",x"1C24");
    gpmc_send('1',x"3395",x"0000");
    gpmc_send('1',x"3396",x"1B25");
    gpmc_send('1',x"3397",x"0000");
    gpmc_send('1',x"3398",x"1A26");
    gpmc_send('1',x"3399",x"0000");
    gpmc_send('1',x"339A",x"1927");
    gpmc_send('1',x"339B",x"0000");
    gpmc_send('1',x"339C",x"1828");
    gpmc_send('1',x"339D",x"0000");
    gpmc_send('1',x"339E",x"1729");
    gpmc_send('1',x"339F",x"0000");
    gpmc_send('1',x"33A0",x"162A");
    gpmc_send('1',x"33A1",x"0000");
    gpmc_send('1',x"33A2",x"152B");
    gpmc_send('1',x"33A3",x"0000");
    gpmc_send('1',x"33A4",x"142C");
    gpmc_send('1',x"33A5",x"0000");
    gpmc_send('1',x"33A6",x"132D");
    gpmc_send('1',x"33A7",x"0000");
    gpmc_send('1',x"33A8",x"122E");
    gpmc_send('1',x"33A9",x"0000");
    gpmc_send('1',x"33AA",x"112F");
    gpmc_send('1',x"33AB",x"0000");
    gpmc_send('1',x"33AC",x"1030");
    gpmc_send('1',x"33AD",x"0000");
    gpmc_send('1',x"33AE",x"0F31");
    gpmc_send('1',x"33AF",x"0000");
    gpmc_send('1',x"33B0",x"0E32");
    gpmc_send('1',x"33B1",x"0000");
    gpmc_send('1',x"33B2",x"0D33");
    gpmc_send('1',x"33B3",x"0000");
    gpmc_send('1',x"33B4",x"0C34");
    gpmc_send('1',x"33B5",x"0000");
    gpmc_send('1',x"33B6",x"0B35");
    gpmc_send('1',x"33B7",x"0000");
    gpmc_send('1',x"33B8",x"0A36");
    gpmc_send('1',x"33B9",x"0000");
    gpmc_send('1',x"33BA",x"0937");
    gpmc_send('1',x"33BB",x"0000");
    gpmc_send('1',x"33BC",x"0838");
    gpmc_send('1',x"33BD",x"0000");
    gpmc_send('1',x"33BE",x"0739");
    gpmc_send('1',x"33BF",x"0000");
    gpmc_send('1',x"33C0",x"063A");
    gpmc_send('1',x"33C1",x"0000");
    gpmc_send('1',x"33C2",x"053B");
    gpmc_send('1',x"33C3",x"0000");
    gpmc_send('1',x"33C4",x"043C");
    gpmc_send('1',x"33C5",x"0000");
    gpmc_send('1',x"33C6",x"033D");
    gpmc_send('1',x"33C7",x"0000");
    gpmc_send('1',x"33C8",x"023E");
    gpmc_send('1',x"33C9",x"0000");
    gpmc_send('1',x"33CA",x"013F");
    gpmc_send('1',x"33CB",x"0000");
    gpmc_send('1',x"33CC",x"003F");
    gpmc_send('1',x"33CD",x"0000");
    gpmc_send('1',x"33CE",x"003E");
    gpmc_send('1',x"33CF",x"0001");
    gpmc_send('1',x"33D0",x"003D");
    gpmc_send('1',x"33D1",x"0002");
    gpmc_send('1',x"33D2",x"003C");
    gpmc_send('1',x"33D3",x"0003");
    gpmc_send('1',x"33D4",x"003B");
    gpmc_send('1',x"33D5",x"0004");
    gpmc_send('1',x"33D6",x"003A");
    gpmc_send('1',x"33D7",x"0005");
    gpmc_send('1',x"33D8",x"0039");
    gpmc_send('1',x"33D9",x"0006");
    gpmc_send('1',x"33DA",x"0038");
    gpmc_send('1',x"33DB",x"0007");
    gpmc_send('1',x"33DC",x"0037");
    gpmc_send('1',x"33DD",x"0008");
    gpmc_send('1',x"33DE",x"0036");
    gpmc_send('1',x"33DF",x"0009");
    gpmc_send('1',x"33E0",x"0035");
    gpmc_send('1',x"33E1",x"000A");
    gpmc_send('1',x"33E2",x"0034");
    gpmc_send('1',x"33E3",x"000B");
    gpmc_send('1',x"33E4",x"0033");
    gpmc_send('1',x"33E5",x"000C");
    gpmc_send('1',x"33E6",x"0032");
    gpmc_send('1',x"33E7",x"000D");
    gpmc_send('1',x"33E8",x"0031");
    gpmc_send('1',x"33E9",x"000E");
    gpmc_send('1',x"33EA",x"0030");
    gpmc_send('1',x"33EB",x"000F");
    gpmc_send('1',x"33EC",x"002F");
    gpmc_send('1',x"33ED",x"0010");
    gpmc_send('1',x"33EE",x"002E");
    gpmc_send('1',x"33EF",x"0011");
    gpmc_send('1',x"33F0",x"002D");
    gpmc_send('1',x"33F1",x"0012");
    gpmc_send('1',x"33F2",x"002C");
    gpmc_send('1',x"33F3",x"0013");
    gpmc_send('1',x"33F4",x"002B");
    gpmc_send('1',x"33F5",x"0014");
    gpmc_send('1',x"33F6",x"002A");
    gpmc_send('1',x"33F7",x"0015");
    gpmc_send('1',x"33F8",x"0029");
    gpmc_send('1',x"33F9",x"0016");
    gpmc_send('1',x"33FA",x"0028");
    gpmc_send('1',x"33FB",x"0017");
    gpmc_send('1',x"33FC",x"0027");
    gpmc_send('1',x"33FD",x"0018");
    gpmc_send('1',x"33FE",x"0026");
    gpmc_send('1',x"33FF",x"0019");
    gpmc_send('1',x"3400",x"0025");
    gpmc_send('1',x"3401",x"001A");
    gpmc_send('1',x"3402",x"0024");
    gpmc_send('1',x"3403",x"001B");
    gpmc_send('1',x"3404",x"0023");
    gpmc_send('1',x"3405",x"001C");
    gpmc_send('1',x"3406",x"0022");
    gpmc_send('1',x"3407",x"001D");
    gpmc_send('1',x"3408",x"0021");
    gpmc_send('1',x"3409",x"001E");
    gpmc_send('1',x"340A",x"0020");
    gpmc_send('1',x"340B",x"001F");
    gpmc_send('1',x"340C",x"001F");
    gpmc_send('1',x"340D",x"0020");
    gpmc_send('1',x"340E",x"001E");
    gpmc_send('1',x"340F",x"0021");
    gpmc_send('1',x"3410",x"001D");
    gpmc_send('1',x"3411",x"0022");
    gpmc_send('1',x"3412",x"001C");
    gpmc_send('1',x"3413",x"0023");
    gpmc_send('1',x"3414",x"001B");
    gpmc_send('1',x"3415",x"0024");
    gpmc_send('1',x"3416",x"001A");
    gpmc_send('1',x"3417",x"0025");
    gpmc_send('1',x"3418",x"0019");
    gpmc_send('1',x"3419",x"0026");
    gpmc_send('1',x"341A",x"0018");
    gpmc_send('1',x"341B",x"0027");
    gpmc_send('1',x"341C",x"0017");
    gpmc_send('1',x"341D",x"0028");
    gpmc_send('1',x"341E",x"0016");
    gpmc_send('1',x"341F",x"0029");
    gpmc_send('1',x"3420",x"0015");
    gpmc_send('1',x"3421",x"002A");
    gpmc_send('1',x"3422",x"0014");
    gpmc_send('1',x"3423",x"002B");
    gpmc_send('1',x"3424",x"0013");
    gpmc_send('1',x"3425",x"002C");
    gpmc_send('1',x"3426",x"0012");
    gpmc_send('1',x"3427",x"002D");
    gpmc_send('1',x"3428",x"0011");
    gpmc_send('1',x"3429",x"002E");
    gpmc_send('1',x"342A",x"0010");
    gpmc_send('1',x"342B",x"002F");
    gpmc_send('1',x"342C",x"000F");
    gpmc_send('1',x"342D",x"0030");
    gpmc_send('1',x"342E",x"000E");
    gpmc_send('1',x"342F",x"0031");
    gpmc_send('1',x"3430",x"000D");
    gpmc_send('1',x"3431",x"0032");
    gpmc_send('1',x"3432",x"000C");
    gpmc_send('1',x"3433",x"0033");
    gpmc_send('1',x"3434",x"000B");
    gpmc_send('1',x"3435",x"0034");
    gpmc_send('1',x"3436",x"000A");
    gpmc_send('1',x"3437",x"0035");
    gpmc_send('1',x"3438",x"0009");
    gpmc_send('1',x"3439",x"0036");
    gpmc_send('1',x"343A",x"0008");
    gpmc_send('1',x"343B",x"0037");
    gpmc_send('1',x"343C",x"0007");
    gpmc_send('1',x"343D",x"0038");
    gpmc_send('1',x"343E",x"0006");
    gpmc_send('1',x"343F",x"0039");
    gpmc_send('1',x"3440",x"0005");
    gpmc_send('1',x"3441",x"003A");
    gpmc_send('1',x"3442",x"0004");
    gpmc_send('1',x"3443",x"003B");
    gpmc_send('1',x"3444",x"0003");
    gpmc_send('1',x"3445",x"003C");
    gpmc_send('1',x"3446",x"0002");
    gpmc_send('1',x"3447",x"003D");
    gpmc_send('1',x"3448",x"0001");
    gpmc_send('1',x"3449",x"003E");
    gpmc_send('1',x"344A",x"0000");
    gpmc_send('1',x"344B",x"003F");
    gpmc_send('1',x"344C",x"0100");
    gpmc_send('1',x"344D",x"003E");
    gpmc_send('1',x"344E",x"0200");
    gpmc_send('1',x"344F",x"003D");
    gpmc_send('1',x"3450",x"0300");
    gpmc_send('1',x"3451",x"003C");
    gpmc_send('1',x"3452",x"0400");
    gpmc_send('1',x"3453",x"003B");
    gpmc_send('1',x"3454",x"0500");
    gpmc_send('1',x"3455",x"003A");
    gpmc_send('1',x"3456",x"0600");
    gpmc_send('1',x"3457",x"0039");
    gpmc_send('1',x"3458",x"0700");
    gpmc_send('1',x"3459",x"0038");
    gpmc_send('1',x"345A",x"0800");
    gpmc_send('1',x"345B",x"0037");
    gpmc_send('1',x"345C",x"0900");
    gpmc_send('1',x"345D",x"0036");
    gpmc_send('1',x"345E",x"0A00");
    gpmc_send('1',x"345F",x"0035");
    gpmc_send('1',x"3460",x"0B00");
    gpmc_send('1',x"3461",x"0034");
    gpmc_send('1',x"3462",x"0C00");
    gpmc_send('1',x"3463",x"0033");
    gpmc_send('1',x"3464",x"0D00");
    gpmc_send('1',x"3465",x"0032");
    gpmc_send('1',x"3466",x"0E00");
    gpmc_send('1',x"3467",x"0031");
    gpmc_send('1',x"3468",x"0F00");
    gpmc_send('1',x"3469",x"0030");
    gpmc_send('1',x"346A",x"1000");
    gpmc_send('1',x"346B",x"002F");
    gpmc_send('1',x"346C",x"1100");
    gpmc_send('1',x"346D",x"002E");
    gpmc_send('1',x"346E",x"1200");
    gpmc_send('1',x"346F",x"002D");
    gpmc_send('1',x"3470",x"1300");
    gpmc_send('1',x"3471",x"002C");
    gpmc_send('1',x"3472",x"1400");
    gpmc_send('1',x"3473",x"002B");
    gpmc_send('1',x"3474",x"1500");
    gpmc_send('1',x"3475",x"002A");
    gpmc_send('1',x"3476",x"1600");
    gpmc_send('1',x"3477",x"0029");
    gpmc_send('1',x"3478",x"1700");
    gpmc_send('1',x"3479",x"0028");
    gpmc_send('1',x"347A",x"1800");
    gpmc_send('1',x"347B",x"0027");
    gpmc_send('1',x"347C",x"1900");
    gpmc_send('1',x"347D",x"0026");
    gpmc_send('1',x"347E",x"1A00");
    gpmc_send('1',x"347F",x"0025");
    gpmc_send('1',x"3480",x"1B00");
    gpmc_send('1',x"3481",x"0024");
    gpmc_send('1',x"3482",x"1C00");
    gpmc_send('1',x"3483",x"0023");
    gpmc_send('1',x"3484",x"1D00");
    gpmc_send('1',x"3485",x"0022");
    gpmc_send('1',x"3486",x"1E00");
    gpmc_send('1',x"3487",x"0021");
    gpmc_send('1',x"3488",x"1F00");
    gpmc_send('1',x"3489",x"0020");
    gpmc_send('1',x"348A",x"2000");
    gpmc_send('1',x"348B",x"001F");
    gpmc_send('1',x"348C",x"2100");
    gpmc_send('1',x"348D",x"001E");
    gpmc_send('1',x"348E",x"2200");
    gpmc_send('1',x"348F",x"001D");
    gpmc_send('1',x"3490",x"2300");
    gpmc_send('1',x"3491",x"001C");
    gpmc_send('1',x"3492",x"2400");
    gpmc_send('1',x"3493",x"001B");
    gpmc_send('1',x"3494",x"2500");
    gpmc_send('1',x"3495",x"001A");
    gpmc_send('1',x"3496",x"2600");
    gpmc_send('1',x"3497",x"0019");
    gpmc_send('1',x"3498",x"2700");
    gpmc_send('1',x"3499",x"0018");
    gpmc_send('1',x"349A",x"2800");
    gpmc_send('1',x"349B",x"0017");
    gpmc_send('1',x"349C",x"2900");
    gpmc_send('1',x"349D",x"0016");
    gpmc_send('1',x"349E",x"2A00");
    gpmc_send('1',x"349F",x"0015");
    gpmc_send('1',x"34A0",x"2B00");
    gpmc_send('1',x"34A1",x"0014");
    gpmc_send('1',x"34A2",x"2C00");
    gpmc_send('1',x"34A3",x"0013");
    gpmc_send('1',x"34A4",x"2D00");
    gpmc_send('1',x"34A5",x"0012");
    gpmc_send('1',x"34A6",x"2E00");
    gpmc_send('1',x"34A7",x"0011");
    gpmc_send('1',x"34A8",x"2F00");
    gpmc_send('1',x"34A9",x"0010");
    gpmc_send('1',x"34AA",x"3000");
    gpmc_send('1',x"34AB",x"000F");
    gpmc_send('1',x"34AC",x"3100");
    gpmc_send('1',x"34AD",x"000E");
    gpmc_send('1',x"34AE",x"3200");
    gpmc_send('1',x"34AF",x"000D");
    gpmc_send('1',x"34B0",x"3300");
    gpmc_send('1',x"34B1",x"000C");
    gpmc_send('1',x"34B2",x"3400");
    gpmc_send('1',x"34B3",x"000B");
    gpmc_send('1',x"34B4",x"3500");
    gpmc_send('1',x"34B5",x"000A");
    gpmc_send('1',x"34B6",x"3600");
    gpmc_send('1',x"34B7",x"0009");
    gpmc_send('1',x"34B8",x"3700");
    gpmc_send('1',x"34B9",x"0008");
    gpmc_send('1',x"34BA",x"3800");
    gpmc_send('1',x"34BB",x"0007");
    gpmc_send('1',x"34BC",x"3900");
    gpmc_send('1',x"34BD",x"0006");
    gpmc_send('1',x"34BE",x"3A00");
    gpmc_send('1',x"34BF",x"0005");
    gpmc_send('1',x"34C0",x"3B00");
    gpmc_send('1',x"34C1",x"0004");
    gpmc_send('1',x"34C2",x"3C00");
    gpmc_send('1',x"34C3",x"0003");
    gpmc_send('1',x"34C4",x"3D00");
    gpmc_send('1',x"34C5",x"0002");
    gpmc_send('1',x"34C6",x"3E00");
    gpmc_send('1',x"34C7",x"0001");
    gpmc_send('1',x"34C8",x"3F00");
    gpmc_send('1',x"34C9",x"0000");
    gpmc_send('1',x"34CA",x"3F01");
    gpmc_send('1',x"34CB",x"0000");
    gpmc_send('1',x"34CC",x"3E02");
    gpmc_send('1',x"34CD",x"0000");
    gpmc_send('1',x"34CE",x"3D03");
    gpmc_send('1',x"34CF",x"0000");
    gpmc_send('1',x"34D0",x"3C04");
    gpmc_send('1',x"34D1",x"0000");
    gpmc_send('1',x"34D2",x"3B05");
    gpmc_send('1',x"34D3",x"0000");
    gpmc_send('1',x"34D4",x"3A06");
    gpmc_send('1',x"34D5",x"0000");
    gpmc_send('1',x"34D6",x"3907");
    gpmc_send('1',x"34D7",x"0000");
    gpmc_send('1',x"34D8",x"3808");
    gpmc_send('1',x"34D9",x"0000");
    gpmc_send('1',x"34DA",x"3709");
    gpmc_send('1',x"34DB",x"0000");
    gpmc_send('1',x"34DC",x"360A");
    gpmc_send('1',x"34DD",x"0000");
    gpmc_send('1',x"34DE",x"350B");
    gpmc_send('1',x"34DF",x"0000");
    gpmc_send('1',x"34E0",x"340C");
    gpmc_send('1',x"34E1",x"0000");
    gpmc_send('1',x"34E2",x"330D");
    gpmc_send('1',x"34E3",x"0000");
    gpmc_send('1',x"34E4",x"320E");
    gpmc_send('1',x"34E5",x"0000");
    gpmc_send('1',x"34E6",x"310F");
    gpmc_send('1',x"34E7",x"0000");
    gpmc_send('1',x"34E8",x"3010");
    gpmc_send('1',x"34E9",x"0000");
    gpmc_send('1',x"34EA",x"2F11");
    gpmc_send('1',x"34EB",x"0000");
    gpmc_send('1',x"34EC",x"2E12");
    gpmc_send('1',x"34ED",x"0000");
    gpmc_send('1',x"34EE",x"2D13");
    gpmc_send('1',x"34EF",x"0000");
    gpmc_send('1',x"34F0",x"2C14");
    gpmc_send('1',x"34F1",x"0000");
    gpmc_send('1',x"34F2",x"2B15");
    gpmc_send('1',x"34F3",x"0000");
    gpmc_send('1',x"34F4",x"2A16");
    gpmc_send('1',x"34F5",x"0000");
    gpmc_send('1',x"34F6",x"2917");
    gpmc_send('1',x"34F7",x"0000");
    gpmc_send('1',x"34F8",x"2818");
    gpmc_send('1',x"34F9",x"0000");
    gpmc_send('1',x"34FA",x"2719");
    gpmc_send('1',x"34FB",x"0000");
    gpmc_send('1',x"34FC",x"261A");
    gpmc_send('1',x"34FD",x"0000");
    gpmc_send('1',x"34FE",x"251B");
    gpmc_send('1',x"34FF",x"0000");
    gpmc_send('1',x"3500",x"241C");
    gpmc_send('1',x"3501",x"0000");
    gpmc_send('1',x"3502",x"231D");
    gpmc_send('1',x"3503",x"0000");
    gpmc_send('1',x"3504",x"221E");
    gpmc_send('1',x"3505",x"0000");
    gpmc_send('1',x"3506",x"211F");
    gpmc_send('1',x"3507",x"0000");
    gpmc_send('1',x"3508",x"2020");
    gpmc_send('1',x"3509",x"0000");
    gpmc_send('1',x"350A",x"1F21");
    gpmc_send('1',x"350B",x"0000");
    gpmc_send('1',x"350C",x"1E22");
    gpmc_send('1',x"350D",x"0000");
    gpmc_send('1',x"350E",x"1D23");
    gpmc_send('1',x"350F",x"0000");
    gpmc_send('1',x"3510",x"1C24");
    gpmc_send('1',x"3511",x"0000");
    gpmc_send('1',x"3512",x"1B25");
    gpmc_send('1',x"3513",x"0000");
    gpmc_send('1',x"3514",x"1A26");
    gpmc_send('1',x"3515",x"0000");
    gpmc_send('1',x"3516",x"1927");
    gpmc_send('1',x"3517",x"0000");
    gpmc_send('1',x"3518",x"1828");
    gpmc_send('1',x"3519",x"0000");
    gpmc_send('1',x"351A",x"1729");
    gpmc_send('1',x"351B",x"0000");
    gpmc_send('1',x"351C",x"162A");
    gpmc_send('1',x"351D",x"0000");
    gpmc_send('1',x"351E",x"152B");
    gpmc_send('1',x"351F",x"0000");
    gpmc_send('1',x"3520",x"142C");
    gpmc_send('1',x"3521",x"0000");
    gpmc_send('1',x"3522",x"132D");
    gpmc_send('1',x"3523",x"0000");
    gpmc_send('1',x"3524",x"122E");
    gpmc_send('1',x"3525",x"0000");
    gpmc_send('1',x"3526",x"112F");
    gpmc_send('1',x"3527",x"0000");
    gpmc_send('1',x"3528",x"1030");
    gpmc_send('1',x"3529",x"0000");
    gpmc_send('1',x"352A",x"0F31");
    gpmc_send('1',x"352B",x"0000");
    gpmc_send('1',x"352C",x"0E32");
    gpmc_send('1',x"352D",x"0000");
    gpmc_send('1',x"352E",x"0D33");
    gpmc_send('1',x"352F",x"0000");
    gpmc_send('1',x"3530",x"0C34");
    gpmc_send('1',x"3531",x"0000");
    gpmc_send('1',x"3532",x"0B35");
    gpmc_send('1',x"3533",x"0000");
    gpmc_send('1',x"3534",x"0A36");
    gpmc_send('1',x"3535",x"0000");
    gpmc_send('1',x"3536",x"0937");
    gpmc_send('1',x"3537",x"0000");
    gpmc_send('1',x"3538",x"0838");
    gpmc_send('1',x"3539",x"0000");
    gpmc_send('1',x"353A",x"0739");
    gpmc_send('1',x"353B",x"0000");
    gpmc_send('1',x"353C",x"063A");
    gpmc_send('1',x"353D",x"0000");
    gpmc_send('1',x"353E",x"053B");
    gpmc_send('1',x"353F",x"0000");
    gpmc_send('1',x"3540",x"043C");
    gpmc_send('1',x"3541",x"0000");
    gpmc_send('1',x"3542",x"033D");
    gpmc_send('1',x"3543",x"0000");
    gpmc_send('1',x"3544",x"023E");
    gpmc_send('1',x"3545",x"0000");
    gpmc_send('1',x"3546",x"013F");
    gpmc_send('1',x"3547",x"0000");
    gpmc_send('1',x"3548",x"003F");
    gpmc_send('1',x"3549",x"0000");
    gpmc_send('1',x"354A",x"003E");
    gpmc_send('1',x"354B",x"0001");
    gpmc_send('1',x"354C",x"003D");
    gpmc_send('1',x"354D",x"0002");
    gpmc_send('1',x"354E",x"003C");
    gpmc_send('1',x"354F",x"0003");
    gpmc_send('1',x"3550",x"003B");
    gpmc_send('1',x"3551",x"0004");
    gpmc_send('1',x"3552",x"003A");
    gpmc_send('1',x"3553",x"0005");
    gpmc_send('1',x"3554",x"0039");
    gpmc_send('1',x"3555",x"0006");
    gpmc_send('1',x"3556",x"0038");
    gpmc_send('1',x"3557",x"0007");
    gpmc_send('1',x"3558",x"0037");
    gpmc_send('1',x"3559",x"0008");
    gpmc_send('1',x"355A",x"0036");
    gpmc_send('1',x"355B",x"0009");
    gpmc_send('1',x"355C",x"0035");
    gpmc_send('1',x"355D",x"000A");
    gpmc_send('1',x"355E",x"0034");
    gpmc_send('1',x"355F",x"000B");
    gpmc_send('1',x"3560",x"0033");
    gpmc_send('1',x"3561",x"000C");
    gpmc_send('1',x"3562",x"0032");
    gpmc_send('1',x"3563",x"000D");
    gpmc_send('1',x"3564",x"0031");
    gpmc_send('1',x"3565",x"000E");
    gpmc_send('1',x"3566",x"0030");
    gpmc_send('1',x"3567",x"000F");
    gpmc_send('1',x"3568",x"002F");
    gpmc_send('1',x"3569",x"0010");
    gpmc_send('1',x"356A",x"002E");
    gpmc_send('1',x"356B",x"0011");
    gpmc_send('1',x"356C",x"002D");
    gpmc_send('1',x"356D",x"0012");
    gpmc_send('1',x"356E",x"002C");
    gpmc_send('1',x"356F",x"0013");
    gpmc_send('1',x"3570",x"002B");
    gpmc_send('1',x"3571",x"0014");
    gpmc_send('1',x"3572",x"002A");
    gpmc_send('1',x"3573",x"0015");
    gpmc_send('1',x"3574",x"0029");
    gpmc_send('1',x"3575",x"0016");
    gpmc_send('1',x"3576",x"0028");
    gpmc_send('1',x"3577",x"0017");
    gpmc_send('1',x"3578",x"0027");
    gpmc_send('1',x"3579",x"0018");
    gpmc_send('1',x"357A",x"0026");
    gpmc_send('1',x"357B",x"0019");
    gpmc_send('1',x"357C",x"0025");
    gpmc_send('1',x"357D",x"001A");
    gpmc_send('1',x"357E",x"0024");
    gpmc_send('1',x"357F",x"001B");
    gpmc_send('1',x"3580",x"0023");
    gpmc_send('1',x"3581",x"001C");
    gpmc_send('1',x"3582",x"0022");
    gpmc_send('1',x"3583",x"001D");
    gpmc_send('1',x"3584",x"0021");
    gpmc_send('1',x"3585",x"001E");
    gpmc_send('1',x"3586",x"0020");
    gpmc_send('1',x"3587",x"001F");
    gpmc_send('1',x"3588",x"001F");
    gpmc_send('1',x"3589",x"0020");
    gpmc_send('1',x"358A",x"001E");
    gpmc_send('1',x"358B",x"0021");
    gpmc_send('1',x"358C",x"001D");
    gpmc_send('1',x"358D",x"0022");
    gpmc_send('1',x"358E",x"001C");
    gpmc_send('1',x"358F",x"0023");
    gpmc_send('1',x"3590",x"001B");
    gpmc_send('1',x"3591",x"0024");
    gpmc_send('1',x"3592",x"001A");
    gpmc_send('1',x"3593",x"0025");
    gpmc_send('1',x"3594",x"0019");
    gpmc_send('1',x"3595",x"0026");
    gpmc_send('1',x"3596",x"0018");
    gpmc_send('1',x"3597",x"0027");
    gpmc_send('1',x"3598",x"0017");
    gpmc_send('1',x"3599",x"0028");
    gpmc_send('1',x"359A",x"0016");
    gpmc_send('1',x"359B",x"0029");
    gpmc_send('1',x"359C",x"0015");
    gpmc_send('1',x"359D",x"002A");
    gpmc_send('1',x"359E",x"0014");
    gpmc_send('1',x"359F",x"002B");
    gpmc_send('1',x"35A0",x"0013");
    gpmc_send('1',x"35A1",x"002C");
    gpmc_send('1',x"35A2",x"0012");
    gpmc_send('1',x"35A3",x"002D");
    gpmc_send('1',x"35A4",x"0011");
    gpmc_send('1',x"35A5",x"002E");
    gpmc_send('1',x"35A6",x"0010");
    gpmc_send('1',x"35A7",x"002F");
    gpmc_send('1',x"35A8",x"000F");
    gpmc_send('1',x"35A9",x"0030");
    gpmc_send('1',x"35AA",x"000E");
    gpmc_send('1',x"35AB",x"0031");
    gpmc_send('1',x"35AC",x"000D");
    gpmc_send('1',x"35AD",x"0032");
    gpmc_send('1',x"35AE",x"000C");
    gpmc_send('1',x"35AF",x"0033");
    gpmc_send('1',x"35B0",x"000B");
    gpmc_send('1',x"35B1",x"0034");
    gpmc_send('1',x"35B2",x"000A");
    gpmc_send('1',x"35B3",x"0035");
    gpmc_send('1',x"35B4",x"0009");
    gpmc_send('1',x"35B5",x"0036");
    gpmc_send('1',x"35B6",x"0008");
    gpmc_send('1',x"35B7",x"0037");
    gpmc_send('1',x"35B8",x"0007");
    gpmc_send('1',x"35B9",x"0038");
    gpmc_send('1',x"35BA",x"0006");
    gpmc_send('1',x"35BB",x"0039");
    gpmc_send('1',x"35BC",x"0005");
    gpmc_send('1',x"35BD",x"003A");
    gpmc_send('1',x"35BE",x"0004");
    gpmc_send('1',x"35BF",x"003B");
    gpmc_send('1',x"35C0",x"0003");
    gpmc_send('1',x"35C1",x"003C");
    gpmc_send('1',x"35C2",x"0002");
    gpmc_send('1',x"35C3",x"003D");
    gpmc_send('1',x"35C4",x"0001");
    gpmc_send('1',x"35C5",x"003E");
    gpmc_send('1',x"35C6",x"0000");
    gpmc_send('1',x"35C7",x"003F");
    gpmc_send('1',x"35C8",x"0100");
    gpmc_send('1',x"35C9",x"003E");
    gpmc_send('1',x"35CA",x"0200");
    gpmc_send('1',x"35CB",x"003D");
    gpmc_send('1',x"35CC",x"0300");
    gpmc_send('1',x"35CD",x"003C");
    gpmc_send('1',x"35CE",x"0400");
    gpmc_send('1',x"35CF",x"003B");
    gpmc_send('1',x"35D0",x"0500");
    gpmc_send('1',x"35D1",x"003A");
    gpmc_send('1',x"35D2",x"0600");
    gpmc_send('1',x"35D3",x"0039");
    gpmc_send('1',x"35D4",x"0700");
    gpmc_send('1',x"35D5",x"0038");
    gpmc_send('1',x"35D6",x"0800");
    gpmc_send('1',x"35D7",x"0037");
    gpmc_send('1',x"35D8",x"0900");
    gpmc_send('1',x"35D9",x"0036");
    gpmc_send('1',x"35DA",x"0A00");
    gpmc_send('1',x"35DB",x"0035");
    gpmc_send('1',x"35DC",x"0B00");
    gpmc_send('1',x"35DD",x"0034");
    gpmc_send('1',x"35DE",x"0C00");
    gpmc_send('1',x"35DF",x"0033");
    gpmc_send('1',x"35E0",x"0D00");
    gpmc_send('1',x"35E1",x"0032");
    gpmc_send('1',x"35E2",x"0E00");
    gpmc_send('1',x"35E3",x"0031");
    gpmc_send('1',x"35E4",x"0F00");
    gpmc_send('1',x"35E5",x"0030");
    gpmc_send('1',x"35E6",x"1000");
    gpmc_send('1',x"35E7",x"002F");
    gpmc_send('1',x"35E8",x"1100");
    gpmc_send('1',x"35E9",x"002E");
    gpmc_send('1',x"35EA",x"1200");
    gpmc_send('1',x"35EB",x"002D");
    gpmc_send('1',x"35EC",x"1300");
    gpmc_send('1',x"35ED",x"002C");
    gpmc_send('1',x"35EE",x"1400");
    gpmc_send('1',x"35EF",x"002B");
    gpmc_send('1',x"35F0",x"1500");
    gpmc_send('1',x"35F1",x"002A");
    gpmc_send('1',x"35F2",x"1600");
    gpmc_send('1',x"35F3",x"0029");
    gpmc_send('1',x"35F4",x"1700");
    gpmc_send('1',x"35F5",x"0028");
    gpmc_send('1',x"35F6",x"1800");
    gpmc_send('1',x"35F7",x"0027");
    gpmc_send('1',x"35F8",x"1900");
    gpmc_send('1',x"35F9",x"0026");
    gpmc_send('1',x"35FA",x"1A00");
    gpmc_send('1',x"35FB",x"0025");
    gpmc_send('1',x"35FC",x"1B00");
    gpmc_send('1',x"35FD",x"0024");
    gpmc_send('1',x"35FE",x"1C00");
    gpmc_send('1',x"35FF",x"0023");
    gpmc_send('1',x"3600",x"1D00");
    gpmc_send('1',x"3601",x"0022");
    gpmc_send('1',x"3602",x"1E00");
    gpmc_send('1',x"3603",x"0021");
    gpmc_send('1',x"3604",x"1F00");
    gpmc_send('1',x"3605",x"0020");
    gpmc_send('1',x"3606",x"2000");
    gpmc_send('1',x"3607",x"001F");
    gpmc_send('1',x"3608",x"2100");
    gpmc_send('1',x"3609",x"001E");
    gpmc_send('1',x"360A",x"2200");
    gpmc_send('1',x"360B",x"001D");
    gpmc_send('1',x"360C",x"2300");
    gpmc_send('1',x"360D",x"001C");
    gpmc_send('1',x"360E",x"2400");
    gpmc_send('1',x"360F",x"001B");
    gpmc_send('1',x"3610",x"2500");
    gpmc_send('1',x"3611",x"001A");
    gpmc_send('1',x"3612",x"2600");
    gpmc_send('1',x"3613",x"0019");
    gpmc_send('1',x"3614",x"2700");
    gpmc_send('1',x"3615",x"0018");
    gpmc_send('1',x"3616",x"2800");
    gpmc_send('1',x"3617",x"0017");
    gpmc_send('1',x"3618",x"2900");
    gpmc_send('1',x"3619",x"0016");
    gpmc_send('1',x"361A",x"2A00");
    gpmc_send('1',x"361B",x"0015");
    gpmc_send('1',x"361C",x"2B00");
    gpmc_send('1',x"361D",x"0014");
    gpmc_send('1',x"361E",x"2C00");
    gpmc_send('1',x"361F",x"0013");
    gpmc_send('1',x"3620",x"2D00");
    gpmc_send('1',x"3621",x"0012");
    gpmc_send('1',x"3622",x"2E00");
    gpmc_send('1',x"3623",x"0011");
    gpmc_send('1',x"3624",x"2F00");
    gpmc_send('1',x"3625",x"0010");
    gpmc_send('1',x"3626",x"3000");
    gpmc_send('1',x"3627",x"000F");
    gpmc_send('1',x"3628",x"3100");
    gpmc_send('1',x"3629",x"000E");
    gpmc_send('1',x"362A",x"3200");
    gpmc_send('1',x"362B",x"000D");
    gpmc_send('1',x"362C",x"3300");
    gpmc_send('1',x"362D",x"000C");
    gpmc_send('1',x"362E",x"3400");
    gpmc_send('1',x"362F",x"000B");
    gpmc_send('1',x"3630",x"3500");
    gpmc_send('1',x"3631",x"000A");
    gpmc_send('1',x"3632",x"3600");
    gpmc_send('1',x"3633",x"0009");
    gpmc_send('1',x"3634",x"3700");
    gpmc_send('1',x"3635",x"0008");
    gpmc_send('1',x"3636",x"3800");
    gpmc_send('1',x"3637",x"0007");
    gpmc_send('1',x"3638",x"3900");
    gpmc_send('1',x"3639",x"0006");
    gpmc_send('1',x"363A",x"3A00");
    gpmc_send('1',x"363B",x"0005");
    gpmc_send('1',x"363C",x"3B00");
    gpmc_send('1',x"363D",x"0004");
    gpmc_send('1',x"363E",x"3C00");
    gpmc_send('1',x"363F",x"0003");
    gpmc_send('1',x"3640",x"3D00");
    gpmc_send('1',x"3641",x"0002");
    gpmc_send('1',x"3642",x"3E00");
    gpmc_send('1',x"3643",x"0001");
    gpmc_send('1',x"3644",x"3F00");
    gpmc_send('1',x"3645",x"0000");
    gpmc_send('1',x"3646",x"3F01");
    gpmc_send('1',x"3647",x"0000");
    gpmc_send('1',x"3648",x"3E02");
    gpmc_send('1',x"3649",x"0000");
    gpmc_send('1',x"364A",x"3D03");
    gpmc_send('1',x"364B",x"0000");
    gpmc_send('1',x"364C",x"3C04");
    gpmc_send('1',x"364D",x"0000");
    gpmc_send('1',x"364E",x"3B05");
    gpmc_send('1',x"364F",x"0000");
    gpmc_send('1',x"3650",x"3A06");
    gpmc_send('1',x"3651",x"0000");
    gpmc_send('1',x"3652",x"3907");
    gpmc_send('1',x"3653",x"0000");
    gpmc_send('1',x"3654",x"3808");
    gpmc_send('1',x"3655",x"0000");
    gpmc_send('1',x"3656",x"3709");
    gpmc_send('1',x"3657",x"0000");
    gpmc_send('1',x"3658",x"360A");
    gpmc_send('1',x"3659",x"0000");
    gpmc_send('1',x"365A",x"350B");
    gpmc_send('1',x"365B",x"0000");
    gpmc_send('1',x"365C",x"340C");
    gpmc_send('1',x"365D",x"0000");
    gpmc_send('1',x"365E",x"330D");
    gpmc_send('1',x"365F",x"0000");
    gpmc_send('1',x"3660",x"320E");
    gpmc_send('1',x"3661",x"0000");
    gpmc_send('1',x"3662",x"310F");
    gpmc_send('1',x"3663",x"0000");
    gpmc_send('1',x"3664",x"3010");
    gpmc_send('1',x"3665",x"0000");
    gpmc_send('1',x"3666",x"2F11");
    gpmc_send('1',x"3667",x"0000");
    gpmc_send('1',x"3668",x"2E12");
    gpmc_send('1',x"3669",x"0000");
    gpmc_send('1',x"366A",x"2D13");
    gpmc_send('1',x"366B",x"0000");
    gpmc_send('1',x"366C",x"2C14");
    gpmc_send('1',x"366D",x"0000");
    gpmc_send('1',x"366E",x"2B15");
    gpmc_send('1',x"366F",x"0000");
    gpmc_send('1',x"3670",x"2A16");
    gpmc_send('1',x"3671",x"0000");
    gpmc_send('1',x"3672",x"2917");
    gpmc_send('1',x"3673",x"0000");
    gpmc_send('1',x"3674",x"2818");
    gpmc_send('1',x"3675",x"0000");
    gpmc_send('1',x"3676",x"2719");
    gpmc_send('1',x"3677",x"0000");
    gpmc_send('1',x"3678",x"261A");
    gpmc_send('1',x"3679",x"0000");
    gpmc_send('1',x"367A",x"251B");
    gpmc_send('1',x"367B",x"0000");
    gpmc_send('1',x"367C",x"241C");
    gpmc_send('1',x"367D",x"0000");
    gpmc_send('1',x"367E",x"231D");
    gpmc_send('1',x"367F",x"0000");
    gpmc_send('1',x"3680",x"221E");
    gpmc_send('1',x"3681",x"0000");
    gpmc_send('1',x"3682",x"211F");
    gpmc_send('1',x"3683",x"0000");
    gpmc_send('1',x"3684",x"2020");
    gpmc_send('1',x"3685",x"0000");
    gpmc_send('1',x"3686",x"1F21");
    gpmc_send('1',x"3687",x"0000");
    gpmc_send('1',x"3688",x"1E22");
    gpmc_send('1',x"3689",x"0000");
    gpmc_send('1',x"368A",x"1D23");
    gpmc_send('1',x"368B",x"0000");
    gpmc_send('1',x"368C",x"1C24");
    gpmc_send('1',x"368D",x"0000");
    gpmc_send('1',x"368E",x"1B25");
    gpmc_send('1',x"368F",x"0000");
    gpmc_send('1',x"3690",x"1A26");
    gpmc_send('1',x"3691",x"0000");
    gpmc_send('1',x"3692",x"1927");
    gpmc_send('1',x"3693",x"0000");
    gpmc_send('1',x"3694",x"1828");
    gpmc_send('1',x"3695",x"0000");
    gpmc_send('1',x"3696",x"1729");
    gpmc_send('1',x"3697",x"0000");
    gpmc_send('1',x"3698",x"162A");
    gpmc_send('1',x"3699",x"0000");
    gpmc_send('1',x"369A",x"152B");
    gpmc_send('1',x"369B",x"0000");
    gpmc_send('1',x"369C",x"142C");
    gpmc_send('1',x"369D",x"0000");
    gpmc_send('1',x"369E",x"132D");
    gpmc_send('1',x"369F",x"0000");
    gpmc_send('1',x"36A0",x"122E");
    gpmc_send('1',x"36A1",x"0000");
    gpmc_send('1',x"36A2",x"112F");
    gpmc_send('1',x"36A3",x"0000");
    gpmc_send('1',x"36A4",x"1030");
    gpmc_send('1',x"36A5",x"0000");
    gpmc_send('1',x"36A6",x"0F31");
    gpmc_send('1',x"36A7",x"0000");
    gpmc_send('1',x"36A8",x"0E32");
    gpmc_send('1',x"36A9",x"0000");
    gpmc_send('1',x"36AA",x"0D33");
    gpmc_send('1',x"36AB",x"0000");
    gpmc_send('1',x"36AC",x"0C34");
    gpmc_send('1',x"36AD",x"0000");
    gpmc_send('1',x"36AE",x"0B35");
    gpmc_send('1',x"36AF",x"0000");
    gpmc_send('1',x"36B0",x"0A36");
    gpmc_send('1',x"36B1",x"0000");
    gpmc_send('1',x"36B2",x"0937");
    gpmc_send('1',x"36B3",x"0000");
    gpmc_send('1',x"36B4",x"0838");
    gpmc_send('1',x"36B5",x"0000");
    gpmc_send('1',x"36B6",x"0739");
    gpmc_send('1',x"36B7",x"0000");
    gpmc_send('1',x"36B8",x"063A");
    gpmc_send('1',x"36B9",x"0000");
    gpmc_send('1',x"36BA",x"053B");
    gpmc_send('1',x"36BB",x"0000");
    gpmc_send('1',x"36BC",x"043C");
    gpmc_send('1',x"36BD",x"0000");
    gpmc_send('1',x"36BE",x"033D");
    gpmc_send('1',x"36BF",x"0000");
    gpmc_send('1',x"36C0",x"023E");
    gpmc_send('1',x"36C1",x"0000");
    gpmc_send('1',x"36C2",x"013F");
    gpmc_send('1',x"36C3",x"0000");
    gpmc_send('1',x"36C4",x"003F");
    gpmc_send('1',x"36C5",x"0000");
    gpmc_send('1',x"36C6",x"003E");
    gpmc_send('1',x"36C7",x"0001");
    gpmc_send('1',x"36C8",x"003D");
    gpmc_send('1',x"36C9",x"0002");
    gpmc_send('1',x"36CA",x"003C");
    gpmc_send('1',x"36CB",x"0003");
    gpmc_send('1',x"36CC",x"003B");
    gpmc_send('1',x"36CD",x"0004");
    gpmc_send('1',x"36CE",x"003A");
    gpmc_send('1',x"36CF",x"0005");
    gpmc_send('1',x"36D0",x"0039");
    gpmc_send('1',x"36D1",x"0006");
    gpmc_send('1',x"36D2",x"0038");
    gpmc_send('1',x"36D3",x"0007");
    gpmc_send('1',x"36D4",x"0037");
    gpmc_send('1',x"36D5",x"0008");
    gpmc_send('1',x"36D6",x"0036");
    gpmc_send('1',x"36D7",x"0009");
    gpmc_send('1',x"36D8",x"0035");
    gpmc_send('1',x"36D9",x"000A");
    gpmc_send('1',x"36DA",x"0034");
    gpmc_send('1',x"36DB",x"000B");
    gpmc_send('1',x"36DC",x"0033");
    gpmc_send('1',x"36DD",x"000C");
    gpmc_send('1',x"36DE",x"0032");
    gpmc_send('1',x"36DF",x"000D");
    gpmc_send('1',x"36E0",x"0031");
    gpmc_send('1',x"36E1",x"000E");
    gpmc_send('1',x"36E2",x"0030");
    gpmc_send('1',x"36E3",x"000F");
    gpmc_send('1',x"36E4",x"002F");
    gpmc_send('1',x"36E5",x"0010");
    gpmc_send('1',x"36E6",x"002E");
    gpmc_send('1',x"36E7",x"0011");
    gpmc_send('1',x"36E8",x"002D");
    gpmc_send('1',x"36E9",x"0012");
    gpmc_send('1',x"36EA",x"002C");
    gpmc_send('1',x"36EB",x"0013");
    gpmc_send('1',x"36EC",x"002B");
    gpmc_send('1',x"36ED",x"0014");
    gpmc_send('1',x"36EE",x"002A");
    gpmc_send('1',x"36EF",x"0015");
    gpmc_send('1',x"36F0",x"0029");
    gpmc_send('1',x"36F1",x"0016");
    gpmc_send('1',x"36F2",x"0028");
    gpmc_send('1',x"36F3",x"0017");
    gpmc_send('1',x"36F4",x"0027");
    gpmc_send('1',x"36F5",x"0018");
    gpmc_send('1',x"36F6",x"0026");
    gpmc_send('1',x"36F7",x"0019");
    gpmc_send('1',x"36F8",x"0025");
    gpmc_send('1',x"36F9",x"001A");
    gpmc_send('1',x"36FA",x"0024");
    gpmc_send('1',x"36FB",x"001B");
    gpmc_send('1',x"36FC",x"0023");
    gpmc_send('1',x"36FD",x"001C");
    gpmc_send('1',x"36FE",x"0022");
    gpmc_send('1',x"36FF",x"001D");
    gpmc_send('1',x"3700",x"0021");
    gpmc_send('1',x"3701",x"001E");
    gpmc_send('1',x"3702",x"0020");
    gpmc_send('1',x"3703",x"001F");
    gpmc_send('1',x"3704",x"001F");
    gpmc_send('1',x"3705",x"0020");
    gpmc_send('1',x"3706",x"001E");
    gpmc_send('1',x"3707",x"0021");
    gpmc_send('1',x"3708",x"001D");
    gpmc_send('1',x"3709",x"0022");
    gpmc_send('1',x"370A",x"001C");
    gpmc_send('1',x"370B",x"0023");
    gpmc_send('1',x"370C",x"001B");
    gpmc_send('1',x"370D",x"0024");
    gpmc_send('1',x"370E",x"001A");
    gpmc_send('1',x"370F",x"0025");
    gpmc_send('1',x"3710",x"0019");
    gpmc_send('1',x"3711",x"0026");
    gpmc_send('1',x"3712",x"0018");
    gpmc_send('1',x"3713",x"0027");
    gpmc_send('1',x"3714",x"0017");
    gpmc_send('1',x"3715",x"0028");
    gpmc_send('1',x"3716",x"0016");
    gpmc_send('1',x"3717",x"0029");
    gpmc_send('1',x"3718",x"0015");
    gpmc_send('1',x"3719",x"002A");
    gpmc_send('1',x"371A",x"0014");
    gpmc_send('1',x"371B",x"002B");
    gpmc_send('1',x"371C",x"0013");
    gpmc_send('1',x"371D",x"002C");
    gpmc_send('1',x"371E",x"0012");
    gpmc_send('1',x"371F",x"002D");
    gpmc_send('1',x"3720",x"0011");
    gpmc_send('1',x"3721",x"002E");
    gpmc_send('1',x"3722",x"0010");
    gpmc_send('1',x"3723",x"002F");
    gpmc_send('1',x"3724",x"000F");
    gpmc_send('1',x"3725",x"0030");
    gpmc_send('1',x"3726",x"000E");
    gpmc_send('1',x"3727",x"0031");
    gpmc_send('1',x"3728",x"000D");
    gpmc_send('1',x"3729",x"0032");
    gpmc_send('1',x"372A",x"000C");
    gpmc_send('1',x"372B",x"0033");
    gpmc_send('1',x"372C",x"000B");
    gpmc_send('1',x"372D",x"0034");
    gpmc_send('1',x"372E",x"000A");
    gpmc_send('1',x"372F",x"0035");
    gpmc_send('1',x"3730",x"0009");
    gpmc_send('1',x"3731",x"0036");
    gpmc_send('1',x"3732",x"0008");
    gpmc_send('1',x"3733",x"0037");
    gpmc_send('1',x"3734",x"0007");
    gpmc_send('1',x"3735",x"0038");
    gpmc_send('1',x"3736",x"0006");
    gpmc_send('1',x"3737",x"0039");
    gpmc_send('1',x"3738",x"0005");
    gpmc_send('1',x"3739",x"003A");
    gpmc_send('1',x"373A",x"0004");
    gpmc_send('1',x"373B",x"003B");
    gpmc_send('1',x"373C",x"0003");
    gpmc_send('1',x"373D",x"003C");
    gpmc_send('1',x"373E",x"0002");
    gpmc_send('1',x"373F",x"003D");
    gpmc_send('1',x"3740",x"0001");
    gpmc_send('1',x"3741",x"003E");
    gpmc_send('1',x"3742",x"0000");
    gpmc_send('1',x"3743",x"003F");
    gpmc_send('1',x"3744",x"0100");
    gpmc_send('1',x"3745",x"003E");
    gpmc_send('1',x"3746",x"0200");
    gpmc_send('1',x"3747",x"003D");
    gpmc_send('1',x"3748",x"0300");
    gpmc_send('1',x"3749",x"003C");
    gpmc_send('1',x"374A",x"0400");
    gpmc_send('1',x"374B",x"003B");
    gpmc_send('1',x"374C",x"0500");
    gpmc_send('1',x"374D",x"003A");
    gpmc_send('1',x"374E",x"0600");
    gpmc_send('1',x"374F",x"0039");
    gpmc_send('1',x"3750",x"0700");
    gpmc_send('1',x"3751",x"0038");
    gpmc_send('1',x"3752",x"0800");
    gpmc_send('1',x"3753",x"0037");
    gpmc_send('1',x"3754",x"0900");
    gpmc_send('1',x"3755",x"0036");
    gpmc_send('1',x"3756",x"0A00");
    gpmc_send('1',x"3757",x"0035");
    gpmc_send('1',x"3758",x"0B00");
    gpmc_send('1',x"3759",x"0034");
    gpmc_send('1',x"375A",x"0C00");
    gpmc_send('1',x"375B",x"0033");
    gpmc_send('1',x"375C",x"0D00");
    gpmc_send('1',x"375D",x"0032");
    gpmc_send('1',x"375E",x"0E00");
    gpmc_send('1',x"375F",x"0031");
    gpmc_send('1',x"3760",x"0F00");
    gpmc_send('1',x"3761",x"0030");
    gpmc_send('1',x"3762",x"1000");
    gpmc_send('1',x"3763",x"002F");
    gpmc_send('1',x"3764",x"1100");
    gpmc_send('1',x"3765",x"002E");
    gpmc_send('1',x"3766",x"1200");
    gpmc_send('1',x"3767",x"002D");
    gpmc_send('1',x"3768",x"1300");
    gpmc_send('1',x"3769",x"002C");
    gpmc_send('1',x"376A",x"1400");
    gpmc_send('1',x"376B",x"002B");
    gpmc_send('1',x"376C",x"1500");
    gpmc_send('1',x"376D",x"002A");
    gpmc_send('1',x"376E",x"1600");
    gpmc_send('1',x"376F",x"0029");
    gpmc_send('1',x"3770",x"1700");
    gpmc_send('1',x"3771",x"0028");
    gpmc_send('1',x"3772",x"1800");
    gpmc_send('1',x"3773",x"0027");
    gpmc_send('1',x"3774",x"1900");
    gpmc_send('1',x"3775",x"0026");
    gpmc_send('1',x"3776",x"1A00");
    gpmc_send('1',x"3777",x"0025");
    gpmc_send('1',x"3778",x"1B00");
    gpmc_send('1',x"3779",x"0024");
    gpmc_send('1',x"377A",x"1C00");
    gpmc_send('1',x"377B",x"0023");
    gpmc_send('1',x"377C",x"1D00");
    gpmc_send('1',x"377D",x"0022");
    gpmc_send('1',x"377E",x"1E00");
    gpmc_send('1',x"377F",x"0021");
    gpmc_send('1',x"3780",x"1F00");
    gpmc_send('1',x"3781",x"0020");
    gpmc_send('1',x"3782",x"2000");
    gpmc_send('1',x"3783",x"001F");
    gpmc_send('1',x"3784",x"2100");
    gpmc_send('1',x"3785",x"001E");
    gpmc_send('1',x"3786",x"2200");
    gpmc_send('1',x"3787",x"001D");
    gpmc_send('1',x"3788",x"2300");
    gpmc_send('1',x"3789",x"001C");
    gpmc_send('1',x"378A",x"2400");
    gpmc_send('1',x"378B",x"001B");
    gpmc_send('1',x"378C",x"2500");
    gpmc_send('1',x"378D",x"001A");
    gpmc_send('1',x"378E",x"2600");
    gpmc_send('1',x"378F",x"0019");
    gpmc_send('1',x"3790",x"2700");
    gpmc_send('1',x"3791",x"0018");
    gpmc_send('1',x"3792",x"2800");
    gpmc_send('1',x"3793",x"0017");
    gpmc_send('1',x"3794",x"2900");
    gpmc_send('1',x"3795",x"0016");
    gpmc_send('1',x"3796",x"2A00");
    gpmc_send('1',x"3797",x"0015");
    gpmc_send('1',x"3798",x"2B00");
    gpmc_send('1',x"3799",x"0014");
    gpmc_send('1',x"379A",x"2C00");
    gpmc_send('1',x"379B",x"0013");
    gpmc_send('1',x"379C",x"2D00");
    gpmc_send('1',x"379D",x"0012");
    gpmc_send('1',x"379E",x"2E00");
    gpmc_send('1',x"379F",x"0011");
    gpmc_send('1',x"37A0",x"2F00");
    gpmc_send('1',x"37A1",x"0010");
    gpmc_send('1',x"37A2",x"3000");
    gpmc_send('1',x"37A3",x"000F");
    gpmc_send('1',x"37A4",x"3100");
    gpmc_send('1',x"37A5",x"000E");
    gpmc_send('1',x"37A6",x"3200");
    gpmc_send('1',x"37A7",x"000D");
    gpmc_send('1',x"37A8",x"3300");
    gpmc_send('1',x"37A9",x"000C");
    gpmc_send('1',x"37AA",x"3400");
    gpmc_send('1',x"37AB",x"000B");
    gpmc_send('1',x"37AC",x"3500");
    gpmc_send('1',x"37AD",x"000A");
    gpmc_send('1',x"37AE",x"3600");
    gpmc_send('1',x"37AF",x"0009");
    gpmc_send('1',x"37B0",x"3700");
    gpmc_send('1',x"37B1",x"0008");
    gpmc_send('1',x"37B2",x"3800");
    gpmc_send('1',x"37B3",x"0007");
    gpmc_send('1',x"37B4",x"3900");
    gpmc_send('1',x"37B5",x"0006");
    gpmc_send('1',x"37B6",x"3A00");
    gpmc_send('1',x"37B7",x"0005");
    gpmc_send('1',x"37B8",x"3B00");
    gpmc_send('1',x"37B9",x"0004");
    gpmc_send('1',x"37BA",x"3C00");
    gpmc_send('1',x"37BB",x"0003");
    gpmc_send('1',x"37BC",x"3D00");
    gpmc_send('1',x"37BD",x"0002");
    gpmc_send('1',x"37BE",x"3E00");
    gpmc_send('1',x"37BF",x"0001");
    gpmc_send('1',x"37C0",x"3F00");
    gpmc_send('1',x"37C1",x"0000");
    gpmc_send('1',x"37C2",x"3F01");
    gpmc_send('1',x"37C3",x"0000");
    gpmc_send('1',x"37C4",x"3E02");
    gpmc_send('1',x"37C5",x"0000");
    gpmc_send('1',x"37C6",x"3D03");
    gpmc_send('1',x"37C7",x"0000");
    gpmc_send('1',x"37C8",x"3C04");
    gpmc_send('1',x"37C9",x"0000");
    gpmc_send('1',x"37CA",x"3B05");
    gpmc_send('1',x"37CB",x"0000");
    gpmc_send('1',x"37CC",x"3A06");
    gpmc_send('1',x"37CD",x"0000");
    gpmc_send('1',x"37CE",x"3907");
    gpmc_send('1',x"37CF",x"0000");
    gpmc_send('1',x"37D0",x"3808");
    gpmc_send('1',x"37D1",x"0000");
    gpmc_send('1',x"37D2",x"3709");
    gpmc_send('1',x"37D3",x"0000");
    gpmc_send('1',x"37D4",x"360A");
    gpmc_send('1',x"37D5",x"0000");
    gpmc_send('1',x"37D6",x"350B");
    gpmc_send('1',x"37D7",x"0000");
    gpmc_send('1',x"37D8",x"340C");
    gpmc_send('1',x"37D9",x"0000");
    gpmc_send('1',x"37DA",x"330D");
    gpmc_send('1',x"37DB",x"0000");
    gpmc_send('1',x"37DC",x"320E");
    gpmc_send('1',x"37DD",x"0000");
    gpmc_send('1',x"37DE",x"310F");
    gpmc_send('1',x"37DF",x"0000");
    gpmc_send('1',x"37E0",x"3010");
    gpmc_send('1',x"37E1",x"0000");
    gpmc_send('1',x"37E2",x"2F11");
    gpmc_send('1',x"37E3",x"0000");
    gpmc_send('1',x"37E4",x"2E12");
    gpmc_send('1',x"37E5",x"0000");
    gpmc_send('1',x"37E6",x"2D13");
    gpmc_send('1',x"37E7",x"0000");
    gpmc_send('1',x"37E8",x"2C14");
    gpmc_send('1',x"37E9",x"0000");
    gpmc_send('1',x"37EA",x"2B15");
    gpmc_send('1',x"37EB",x"0000");
    gpmc_send('1',x"37EC",x"2A16");
    gpmc_send('1',x"37ED",x"0000");
    gpmc_send('1',x"37EE",x"2917");
    gpmc_send('1',x"37EF",x"0000");
    gpmc_send('1',x"37F0",x"2818");
    gpmc_send('1',x"37F1",x"0000");
    gpmc_send('1',x"37F2",x"2719");
    gpmc_send('1',x"37F3",x"0000");
    gpmc_send('1',x"37F4",x"261A");
    gpmc_send('1',x"37F5",x"0000");
    gpmc_send('1',x"37F6",x"251B");
    gpmc_send('1',x"37F7",x"0000");
    gpmc_send('1',x"37F8",x"241C");
    gpmc_send('1',x"37F9",x"0000");
    gpmc_send('1',x"37FA",x"231D");
    gpmc_send('1',x"37FB",x"0000");
    gpmc_send('1',x"37FC",x"221E");
    gpmc_send('1',x"37FD",x"0000");
    gpmc_send('1',x"37FE",x"211F");
    gpmc_send('1',x"37FF",x"0000");
    gpmc_send('1',x"3800",x"2020");
    gpmc_send('1',x"3801",x"0000");
    gpmc_send('1',x"3802",x"1F21");
    gpmc_send('1',x"3803",x"0000");
    gpmc_send('1',x"3804",x"1E22");
    gpmc_send('1',x"3805",x"0000");
    gpmc_send('1',x"3806",x"1D23");
    gpmc_send('1',x"3807",x"0000");
    gpmc_send('1',x"3808",x"1C24");
    gpmc_send('1',x"3809",x"0000");
    gpmc_send('1',x"380A",x"1B25");
    gpmc_send('1',x"380B",x"0000");
    gpmc_send('1',x"380C",x"1A26");
    gpmc_send('1',x"380D",x"0000");
    gpmc_send('1',x"380E",x"1927");
    gpmc_send('1',x"380F",x"0000");
    gpmc_send('1',x"3810",x"1828");
    gpmc_send('1',x"3811",x"0000");
    gpmc_send('1',x"3812",x"1729");
    gpmc_send('1',x"3813",x"0000");
    gpmc_send('1',x"3814",x"162A");
    gpmc_send('1',x"3815",x"0000");
    gpmc_send('1',x"3816",x"152B");
    gpmc_send('1',x"3817",x"0000");
    gpmc_send('1',x"3818",x"142C");
    gpmc_send('1',x"3819",x"0000");
    gpmc_send('1',x"381A",x"132D");
    gpmc_send('1',x"381B",x"0000");
    gpmc_send('1',x"381C",x"122E");
    gpmc_send('1',x"381D",x"0000");
    gpmc_send('1',x"381E",x"112F");
    gpmc_send('1',x"381F",x"0000");
    gpmc_send('1',x"3820",x"1030");
    gpmc_send('1',x"3821",x"0000");
    gpmc_send('1',x"3822",x"0F31");
    gpmc_send('1',x"3823",x"0000");
    gpmc_send('1',x"3824",x"0E32");
    gpmc_send('1',x"3825",x"0000");
    gpmc_send('1',x"3826",x"0D33");
    gpmc_send('1',x"3827",x"0000");
    gpmc_send('1',x"3828",x"0C34");
    gpmc_send('1',x"3829",x"0000");
    gpmc_send('1',x"382A",x"0B35");
    gpmc_send('1',x"382B",x"0000");
    gpmc_send('1',x"382C",x"0A36");
    gpmc_send('1',x"382D",x"0000");
    gpmc_send('1',x"382E",x"0937");
    gpmc_send('1',x"382F",x"0000");
    gpmc_send('1',x"3830",x"0838");
    gpmc_send('1',x"3831",x"0000");
    gpmc_send('1',x"3832",x"0739");
    gpmc_send('1',x"3833",x"0000");
    gpmc_send('1',x"3834",x"063A");
    gpmc_send('1',x"3835",x"0000");
    gpmc_send('1',x"3836",x"053B");
    gpmc_send('1',x"3837",x"0000");
    gpmc_send('1',x"3838",x"043C");
    gpmc_send('1',x"3839",x"0000");
    gpmc_send('1',x"383A",x"033D");
    gpmc_send('1',x"383B",x"0000");
    gpmc_send('1',x"383C",x"023E");
    gpmc_send('1',x"383D",x"0000");
    gpmc_send('1',x"383E",x"013F");
    gpmc_send('1',x"383F",x"0000");
    gpmc_send('1',x"3840",x"003F");
    gpmc_send('1',x"3841",x"0000");
    gpmc_send('1',x"3842",x"003E");
    gpmc_send('1',x"3843",x"0001");
    gpmc_send('1',x"3844",x"003D");
    gpmc_send('1',x"3845",x"0002");
    gpmc_send('1',x"3846",x"003C");
    gpmc_send('1',x"3847",x"0003");
    gpmc_send('1',x"3848",x"003B");
    gpmc_send('1',x"3849",x"0004");
    gpmc_send('1',x"384A",x"003A");
    gpmc_send('1',x"384B",x"0005");
    gpmc_send('1',x"384C",x"0039");
    gpmc_send('1',x"384D",x"0006");
    gpmc_send('1',x"384E",x"0038");
    gpmc_send('1',x"384F",x"0007");
    gpmc_send('1',x"3850",x"0037");
    gpmc_send('1',x"3851",x"0008");
    gpmc_send('1',x"3852",x"0036");
    gpmc_send('1',x"3853",x"0009");
    gpmc_send('1',x"3854",x"0035");
    gpmc_send('1',x"3855",x"000A");
    gpmc_send('1',x"3856",x"0034");
    gpmc_send('1',x"3857",x"000B");
    gpmc_send('1',x"3858",x"0033");
    gpmc_send('1',x"3859",x"000C");
    gpmc_send('1',x"385A",x"0032");
    gpmc_send('1',x"385B",x"000D");
    gpmc_send('1',x"385C",x"0031");
    gpmc_send('1',x"385D",x"000E");
    gpmc_send('1',x"385E",x"0030");
    gpmc_send('1',x"385F",x"000F");
    gpmc_send('1',x"3860",x"002F");
    gpmc_send('1',x"3861",x"0010");
    gpmc_send('1',x"3862",x"002E");
    gpmc_send('1',x"3863",x"0011");
    gpmc_send('1',x"3864",x"002D");
    gpmc_send('1',x"3865",x"0012");
    gpmc_send('1',x"3866",x"002C");
    gpmc_send('1',x"3867",x"0013");
    gpmc_send('1',x"3868",x"002B");
    gpmc_send('1',x"3869",x"0014");
    gpmc_send('1',x"386A",x"002A");
    gpmc_send('1',x"386B",x"0015");
    gpmc_send('1',x"386C",x"0029");
    gpmc_send('1',x"386D",x"0016");
    gpmc_send('1',x"386E",x"0028");
    gpmc_send('1',x"386F",x"0017");
    gpmc_send('1',x"3870",x"0027");
    gpmc_send('1',x"3871",x"0018");
    gpmc_send('1',x"3872",x"0026");
    gpmc_send('1',x"3873",x"0019");
    gpmc_send('1',x"3874",x"0025");
    gpmc_send('1',x"3875",x"001A");
    gpmc_send('1',x"3876",x"0024");
    gpmc_send('1',x"3877",x"001B");
    gpmc_send('1',x"3878",x"0023");
    gpmc_send('1',x"3879",x"001C");
    gpmc_send('1',x"387A",x"0022");
    gpmc_send('1',x"387B",x"001D");
    gpmc_send('1',x"387C",x"0021");
    gpmc_send('1',x"387D",x"001E");
    gpmc_send('1',x"387E",x"0020");
    gpmc_send('1',x"387F",x"001F");
    gpmc_send('1',x"3880",x"001F");
    gpmc_send('1',x"3881",x"0020");
    gpmc_send('1',x"3882",x"001E");
    gpmc_send('1',x"3883",x"0021");
    gpmc_send('1',x"3884",x"001D");
    gpmc_send('1',x"3885",x"0022");
    gpmc_send('1',x"3886",x"001C");
    gpmc_send('1',x"3887",x"0023");
    gpmc_send('1',x"3888",x"001B");
    gpmc_send('1',x"3889",x"0024");
    gpmc_send('1',x"388A",x"001A");
    gpmc_send('1',x"388B",x"0025");
    gpmc_send('1',x"388C",x"0019");
    gpmc_send('1',x"388D",x"0026");
    gpmc_send('1',x"388E",x"0018");
    gpmc_send('1',x"388F",x"0027");
    gpmc_send('1',x"3890",x"0017");
    gpmc_send('1',x"3891",x"0028");
    gpmc_send('1',x"3892",x"0016");
    gpmc_send('1',x"3893",x"0029");
    gpmc_send('1',x"3894",x"0015");
    gpmc_send('1',x"3895",x"002A");
    gpmc_send('1',x"3896",x"0014");
    gpmc_send('1',x"3897",x"002B");
    gpmc_send('1',x"3898",x"0013");
    gpmc_send('1',x"3899",x"002C");
    gpmc_send('1',x"389A",x"0012");
    gpmc_send('1',x"389B",x"002D");
    gpmc_send('1',x"389C",x"0011");
    gpmc_send('1',x"389D",x"002E");
    gpmc_send('1',x"389E",x"0010");
    gpmc_send('1',x"389F",x"002F");
    gpmc_send('1',x"38A0",x"000F");
    gpmc_send('1',x"38A1",x"0030");
    gpmc_send('1',x"38A2",x"000E");
    gpmc_send('1',x"38A3",x"0031");
    gpmc_send('1',x"38A4",x"000D");
    gpmc_send('1',x"38A5",x"0032");
    gpmc_send('1',x"38A6",x"000C");
    gpmc_send('1',x"38A7",x"0033");
    gpmc_send('1',x"38A8",x"000B");
    gpmc_send('1',x"38A9",x"0034");
    gpmc_send('1',x"38AA",x"000A");
    gpmc_send('1',x"38AB",x"0035");
    gpmc_send('1',x"38AC",x"0009");
    gpmc_send('1',x"38AD",x"0036");
    gpmc_send('1',x"38AE",x"0008");
    gpmc_send('1',x"38AF",x"0037");
    gpmc_send('1',x"38B0",x"0007");
    gpmc_send('1',x"38B1",x"0038");
    gpmc_send('1',x"38B2",x"0006");
    gpmc_send('1',x"38B3",x"0039");
    gpmc_send('1',x"38B4",x"0005");
    gpmc_send('1',x"38B5",x"003A");
    gpmc_send('1',x"38B6",x"0004");
    gpmc_send('1',x"38B7",x"003B");
    gpmc_send('1',x"38B8",x"0003");
    gpmc_send('1',x"38B9",x"003C");
    gpmc_send('1',x"38BA",x"0002");
    gpmc_send('1',x"38BB",x"003D");
    gpmc_send('1',x"38BC",x"0001");
    gpmc_send('1',x"38BD",x"003E");
    gpmc_send('1',x"38BE",x"0000");
    gpmc_send('1',x"38BF",x"003F");
    gpmc_send('1',x"38C0",x"0100");
    gpmc_send('1',x"38C1",x"003E");
    gpmc_send('1',x"38C2",x"0200");
    gpmc_send('1',x"38C3",x"003D");
    gpmc_send('1',x"38C4",x"0300");
    gpmc_send('1',x"38C5",x"003C");
    gpmc_send('1',x"38C6",x"0400");
    gpmc_send('1',x"38C7",x"003B");
    gpmc_send('1',x"38C8",x"0500");
    gpmc_send('1',x"38C9",x"003A");
    gpmc_send('1',x"38CA",x"0600");
    gpmc_send('1',x"38CB",x"0039");
    gpmc_send('1',x"38CC",x"0700");
    gpmc_send('1',x"38CD",x"0038");
    gpmc_send('1',x"38CE",x"0800");
    gpmc_send('1',x"38CF",x"0037");
    gpmc_send('1',x"38D0",x"0900");
    gpmc_send('1',x"38D1",x"0036");
    gpmc_send('1',x"38D2",x"0A00");
    gpmc_send('1',x"38D3",x"0035");
    gpmc_send('1',x"38D4",x"0B00");
    gpmc_send('1',x"38D5",x"0034");
    gpmc_send('1',x"38D6",x"0C00");
    gpmc_send('1',x"38D7",x"0033");
    gpmc_send('1',x"38D8",x"0D00");
    gpmc_send('1',x"38D9",x"0032");
    gpmc_send('1',x"38DA",x"0E00");
    gpmc_send('1',x"38DB",x"0031");
    gpmc_send('1',x"38DC",x"0F00");
    gpmc_send('1',x"38DD",x"0030");
    gpmc_send('1',x"38DE",x"1000");
    gpmc_send('1',x"38DF",x"002F");
    gpmc_send('1',x"38E0",x"1100");
    gpmc_send('1',x"38E1",x"002E");
    gpmc_send('1',x"38E2",x"1200");
    gpmc_send('1',x"38E3",x"002D");
    gpmc_send('1',x"38E4",x"1300");
    gpmc_send('1',x"38E5",x"002C");
    gpmc_send('1',x"38E6",x"1400");
    gpmc_send('1',x"38E7",x"002B");
    gpmc_send('1',x"38E8",x"1500");
    gpmc_send('1',x"38E9",x"002A");
    gpmc_send('1',x"38EA",x"1600");
    gpmc_send('1',x"38EB",x"0029");
    gpmc_send('1',x"38EC",x"1700");
    gpmc_send('1',x"38ED",x"0028");
    gpmc_send('1',x"38EE",x"1800");
    gpmc_send('1',x"38EF",x"0027");
    gpmc_send('1',x"38F0",x"1900");
    gpmc_send('1',x"38F1",x"0026");
    gpmc_send('1',x"38F2",x"1A00");
    gpmc_send('1',x"38F3",x"0025");
    gpmc_send('1',x"38F4",x"1B00");
    gpmc_send('1',x"38F5",x"0024");
    gpmc_send('1',x"38F6",x"1C00");
    gpmc_send('1',x"38F7",x"0023");
    gpmc_send('1',x"38F8",x"1D00");
    gpmc_send('1',x"38F9",x"0022");
    gpmc_send('1',x"38FA",x"1E00");
    gpmc_send('1',x"38FB",x"0021");
    gpmc_send('1',x"38FC",x"1F00");
    gpmc_send('1',x"38FD",x"0020");
    gpmc_send('1',x"38FE",x"2000");
    gpmc_send('1',x"38FF",x"001F");
    gpmc_send('1',x"3900",x"2100");
    gpmc_send('1',x"3901",x"001E");
    gpmc_send('1',x"3902",x"2200");
    gpmc_send('1',x"3903",x"001D");
    gpmc_send('1',x"3904",x"2300");
    gpmc_send('1',x"3905",x"001C");
    gpmc_send('1',x"3906",x"2400");
    gpmc_send('1',x"3907",x"001B");
    gpmc_send('1',x"3908",x"2500");
    gpmc_send('1',x"3909",x"001A");
    gpmc_send('1',x"390A",x"2600");
    gpmc_send('1',x"390B",x"0019");
    gpmc_send('1',x"390C",x"2700");
    gpmc_send('1',x"390D",x"0018");
    gpmc_send('1',x"390E",x"2800");
    gpmc_send('1',x"390F",x"0017");
    gpmc_send('1',x"3910",x"2900");
    gpmc_send('1',x"3911",x"0016");
    gpmc_send('1',x"3912",x"2A00");
    gpmc_send('1',x"3913",x"0015");
    gpmc_send('1',x"3914",x"2B00");
    gpmc_send('1',x"3915",x"0014");
    gpmc_send('1',x"3916",x"2C00");
    gpmc_send('1',x"3917",x"0013");
    gpmc_send('1',x"3918",x"2D00");
    gpmc_send('1',x"3919",x"0012");
    gpmc_send('1',x"391A",x"2E00");
    gpmc_send('1',x"391B",x"0011");
    gpmc_send('1',x"391C",x"2F00");
    gpmc_send('1',x"391D",x"0010");
    gpmc_send('1',x"391E",x"3000");
    gpmc_send('1',x"391F",x"000F");
    gpmc_send('1',x"3920",x"3100");
    gpmc_send('1',x"3921",x"000E");
    gpmc_send('1',x"3922",x"3200");
    gpmc_send('1',x"3923",x"000D");
    gpmc_send('1',x"3924",x"3300");
    gpmc_send('1',x"3925",x"000C");
    gpmc_send('1',x"3926",x"3400");
    gpmc_send('1',x"3927",x"000B");
    gpmc_send('1',x"3928",x"3500");
    gpmc_send('1',x"3929",x"000A");
    gpmc_send('1',x"392A",x"3600");
    gpmc_send('1',x"392B",x"0009");
    gpmc_send('1',x"392C",x"3700");
    gpmc_send('1',x"392D",x"0008");
    gpmc_send('1',x"392E",x"3800");
    gpmc_send('1',x"392F",x"0007");
    gpmc_send('1',x"3930",x"3900");
    gpmc_send('1',x"3931",x"0006");
    gpmc_send('1',x"3932",x"3A00");
    gpmc_send('1',x"3933",x"0005");
    gpmc_send('1',x"3934",x"3B00");
    gpmc_send('1',x"3935",x"0004");
    gpmc_send('1',x"3936",x"3C00");
    gpmc_send('1',x"3937",x"0003");
    gpmc_send('1',x"3938",x"3D00");
    gpmc_send('1',x"3939",x"0002");
    gpmc_send('1',x"393A",x"3E00");
    gpmc_send('1',x"393B",x"0001");
    gpmc_send('1',x"393C",x"3F00");
    gpmc_send('1',x"393D",x"0000");
    gpmc_send('1',x"393E",x"3F01");
    gpmc_send('1',x"393F",x"0000");
    gpmc_send('1',x"3940",x"3E02");
    gpmc_send('1',x"3941",x"0000");
    gpmc_send('1',x"3942",x"3D03");
    gpmc_send('1',x"3943",x"0000");
    gpmc_send('1',x"3944",x"3C04");
    gpmc_send('1',x"3945",x"0000");
    gpmc_send('1',x"3946",x"3B05");
    gpmc_send('1',x"3947",x"0000");
    gpmc_send('1',x"3948",x"3A06");
    gpmc_send('1',x"3949",x"0000");
    gpmc_send('1',x"394A",x"3907");
    gpmc_send('1',x"394B",x"0000");
    gpmc_send('1',x"394C",x"3808");
    gpmc_send('1',x"394D",x"0000");
    gpmc_send('1',x"394E",x"3709");
    gpmc_send('1',x"394F",x"0000");
    gpmc_send('1',x"3950",x"360A");
    gpmc_send('1',x"3951",x"0000");
    gpmc_send('1',x"3952",x"350B");
    gpmc_send('1',x"3953",x"0000");
    gpmc_send('1',x"3954",x"340C");
    gpmc_send('1',x"3955",x"0000");
    gpmc_send('1',x"3956",x"330D");
    gpmc_send('1',x"3957",x"0000");
    gpmc_send('1',x"3958",x"320E");
    gpmc_send('1',x"3959",x"0000");
    gpmc_send('1',x"395A",x"310F");
    gpmc_send('1',x"395B",x"0000");
    gpmc_send('1',x"395C",x"3010");
    gpmc_send('1',x"395D",x"0000");
    gpmc_send('1',x"395E",x"2F11");
    gpmc_send('1',x"395F",x"0000");
    gpmc_send('1',x"3960",x"2E12");
    gpmc_send('1',x"3961",x"0000");
    gpmc_send('1',x"3962",x"2D13");
    gpmc_send('1',x"3963",x"0000");
    gpmc_send('1',x"3964",x"2C14");
    gpmc_send('1',x"3965",x"0000");
    gpmc_send('1',x"3966",x"2B15");
    gpmc_send('1',x"3967",x"0000");
    gpmc_send('1',x"3968",x"2A16");
    gpmc_send('1',x"3969",x"0000");
    gpmc_send('1',x"396A",x"2917");
    gpmc_send('1',x"396B",x"0000");
    gpmc_send('1',x"396C",x"2818");
    gpmc_send('1',x"396D",x"0000");
    gpmc_send('1',x"396E",x"2719");
    gpmc_send('1',x"396F",x"0000");
    gpmc_send('1',x"3970",x"261A");
    gpmc_send('1',x"3971",x"0000");
    gpmc_send('1',x"3972",x"251B");
    gpmc_send('1',x"3973",x"0000");
    gpmc_send('1',x"3974",x"241C");
    gpmc_send('1',x"3975",x"0000");
    gpmc_send('1',x"3976",x"231D");
    gpmc_send('1',x"3977",x"0000");
    gpmc_send('1',x"3978",x"221E");
    gpmc_send('1',x"3979",x"0000");
    gpmc_send('1',x"397A",x"211F");
    gpmc_send('1',x"397B",x"0000");
    gpmc_send('1',x"397C",x"2020");
    gpmc_send('1',x"397D",x"0000");
    gpmc_send('1',x"397E",x"1F21");
    gpmc_send('1',x"397F",x"0000");
    gpmc_send('1',x"3980",x"1E22");
    gpmc_send('1',x"3981",x"0000");
    gpmc_send('1',x"3982",x"1D23");
    gpmc_send('1',x"3983",x"0000");
    gpmc_send('1',x"3984",x"1C24");
    gpmc_send('1',x"3985",x"0000");
    gpmc_send('1',x"3986",x"1B25");
    gpmc_send('1',x"3987",x"0000");
    gpmc_send('1',x"3988",x"1A26");
    gpmc_send('1',x"3989",x"0000");
    gpmc_send('1',x"398A",x"1927");
    gpmc_send('1',x"398B",x"0000");
    gpmc_send('1',x"398C",x"1828");
    gpmc_send('1',x"398D",x"0000");
    gpmc_send('1',x"398E",x"1729");
    gpmc_send('1',x"398F",x"0000");
    gpmc_send('1',x"3990",x"162A");
    gpmc_send('1',x"3991",x"0000");
    gpmc_send('1',x"3992",x"152B");
    gpmc_send('1',x"3993",x"0000");
    gpmc_send('1',x"3994",x"142C");
    gpmc_send('1',x"3995",x"0000");
    gpmc_send('1',x"3996",x"132D");
    gpmc_send('1',x"3997",x"0000");
    gpmc_send('1',x"3998",x"122E");
    gpmc_send('1',x"3999",x"0000");
    gpmc_send('1',x"399A",x"112F");
    gpmc_send('1',x"399B",x"0000");
    gpmc_send('1',x"399C",x"1030");
    gpmc_send('1',x"399D",x"0000");
    gpmc_send('1',x"399E",x"0F31");
    gpmc_send('1',x"399F",x"0000");
    gpmc_send('1',x"39A0",x"0E32");
    gpmc_send('1',x"39A1",x"0000");
    gpmc_send('1',x"39A2",x"0D33");
    gpmc_send('1',x"39A3",x"0000");
    gpmc_send('1',x"39A4",x"0C34");
    gpmc_send('1',x"39A5",x"0000");
    gpmc_send('1',x"39A6",x"0B35");
    gpmc_send('1',x"39A7",x"0000");
    gpmc_send('1',x"39A8",x"0A36");
    gpmc_send('1',x"39A9",x"0000");
    gpmc_send('1',x"39AA",x"0937");
    gpmc_send('1',x"39AB",x"0000");
    gpmc_send('1',x"39AC",x"0838");
    gpmc_send('1',x"39AD",x"0000");
    gpmc_send('1',x"39AE",x"0739");
    gpmc_send('1',x"39AF",x"0000");
    gpmc_send('1',x"39B0",x"063A");
    gpmc_send('1',x"39B1",x"0000");
    gpmc_send('1',x"39B2",x"053B");
    gpmc_send('1',x"39B3",x"0000");
    gpmc_send('1',x"39B4",x"043C");
    gpmc_send('1',x"39B5",x"0000");
    gpmc_send('1',x"39B6",x"033D");
    gpmc_send('1',x"39B7",x"0000");
    gpmc_send('1',x"39B8",x"023E");
    gpmc_send('1',x"39B9",x"0000");
    gpmc_send('1',x"39BA",x"013F");
    gpmc_send('1',x"39BB",x"0000");
    gpmc_send('1',x"39BC",x"003F");
    gpmc_send('1',x"39BD",x"0000");
    gpmc_send('1',x"39BE",x"003E");
    gpmc_send('1',x"39BF",x"0001");
    gpmc_send('1',x"39C0",x"003D");
    gpmc_send('1',x"39C1",x"0002");
    gpmc_send('1',x"39C2",x"003C");
    gpmc_send('1',x"39C3",x"0003");
    gpmc_send('1',x"39C4",x"003B");
    gpmc_send('1',x"39C5",x"0004");
    gpmc_send('1',x"39C6",x"003A");
    gpmc_send('1',x"39C7",x"0005");
    gpmc_send('1',x"39C8",x"0039");
    gpmc_send('1',x"39C9",x"0006");
    gpmc_send('1',x"39CA",x"0038");
    gpmc_send('1',x"39CB",x"0007");
    gpmc_send('1',x"39CC",x"0037");
    gpmc_send('1',x"39CD",x"0008");
    gpmc_send('1',x"39CE",x"0036");
    gpmc_send('1',x"39CF",x"0009");
    gpmc_send('1',x"39D0",x"0035");
    gpmc_send('1',x"39D1",x"000A");
    gpmc_send('1',x"39D2",x"0034");
    gpmc_send('1',x"39D3",x"000B");
    gpmc_send('1',x"39D4",x"0033");
    gpmc_send('1',x"39D5",x"000C");
    gpmc_send('1',x"39D6",x"0032");
    gpmc_send('1',x"39D7",x"000D");
    gpmc_send('1',x"39D8",x"0031");
    gpmc_send('1',x"39D9",x"000E");
    gpmc_send('1',x"39DA",x"0030");
    gpmc_send('1',x"39DB",x"000F");
    gpmc_send('1',x"39DC",x"002F");
    gpmc_send('1',x"39DD",x"0010");
    gpmc_send('1',x"39DE",x"002E");
    gpmc_send('1',x"39DF",x"0011");
    gpmc_send('1',x"39E0",x"002D");
    gpmc_send('1',x"39E1",x"0012");
    gpmc_send('1',x"39E2",x"002C");
    gpmc_send('1',x"39E3",x"0013");
    gpmc_send('1',x"39E4",x"002B");
    gpmc_send('1',x"39E5",x"0014");
    gpmc_send('1',x"39E6",x"002A");
    gpmc_send('1',x"39E7",x"0015");
    gpmc_send('1',x"39E8",x"0029");
    gpmc_send('1',x"39E9",x"0016");
    gpmc_send('1',x"39EA",x"0028");
    gpmc_send('1',x"39EB",x"0017");
    gpmc_send('1',x"39EC",x"0027");
    gpmc_send('1',x"39ED",x"0018");
    gpmc_send('1',x"39EE",x"0026");
    gpmc_send('1',x"39EF",x"0019");
    gpmc_send('1',x"39F0",x"0025");
    gpmc_send('1',x"39F1",x"001A");
    gpmc_send('1',x"39F2",x"0024");
    gpmc_send('1',x"39F3",x"001B");
    gpmc_send('1',x"39F4",x"0023");
    gpmc_send('1',x"39F5",x"001C");
    gpmc_send('1',x"39F6",x"0022");
    gpmc_send('1',x"39F7",x"001D");
    gpmc_send('1',x"39F8",x"0021");
    gpmc_send('1',x"39F9",x"001E");
    gpmc_send('1',x"39FA",x"0020");
    gpmc_send('1',x"39FB",x"001F");
    gpmc_send('1',x"39FC",x"001F");
    gpmc_send('1',x"39FD",x"0020");
    gpmc_send('1',x"39FE",x"001E");
    gpmc_send('1',x"39FF",x"0021");
    gpmc_send('1',x"3A00",x"001D");
    gpmc_send('1',x"3A01",x"0022");
    gpmc_send('1',x"3A02",x"001C");
    gpmc_send('1',x"3A03",x"0023");
    gpmc_send('1',x"3A04",x"001B");
    gpmc_send('1',x"3A05",x"0024");
    gpmc_send('1',x"3A06",x"001A");
    gpmc_send('1',x"3A07",x"0025");
    gpmc_send('1',x"3A08",x"0019");
    gpmc_send('1',x"3A09",x"0026");
    gpmc_send('1',x"3A0A",x"0018");
    gpmc_send('1',x"3A0B",x"0027");
    gpmc_send('1',x"3A0C",x"0017");
    gpmc_send('1',x"3A0D",x"0028");
    gpmc_send('1',x"3A0E",x"0016");
    gpmc_send('1',x"3A0F",x"0029");
    gpmc_send('1',x"3A10",x"0015");
    gpmc_send('1',x"3A11",x"002A");
    gpmc_send('1',x"3A12",x"0014");
    gpmc_send('1',x"3A13",x"002B");
    gpmc_send('1',x"3A14",x"0013");
    gpmc_send('1',x"3A15",x"002C");
    gpmc_send('1',x"3A16",x"0012");
    gpmc_send('1',x"3A17",x"002D");
    gpmc_send('1',x"3A18",x"0011");
    gpmc_send('1',x"3A19",x"002E");
    gpmc_send('1',x"3A1A",x"0010");
    gpmc_send('1',x"3A1B",x"002F");
    gpmc_send('1',x"3A1C",x"000F");
    gpmc_send('1',x"3A1D",x"0030");
    gpmc_send('1',x"3A1E",x"000E");
    gpmc_send('1',x"3A1F",x"0031");
    gpmc_send('1',x"3A20",x"000D");
    gpmc_send('1',x"3A21",x"0032");
    gpmc_send('1',x"3A22",x"000C");
    gpmc_send('1',x"3A23",x"0033");
    gpmc_send('1',x"3A24",x"000B");
    gpmc_send('1',x"3A25",x"0034");
    gpmc_send('1',x"3A26",x"000A");
    gpmc_send('1',x"3A27",x"0035");
    gpmc_send('1',x"3A28",x"0009");
    gpmc_send('1',x"3A29",x"0036");
    gpmc_send('1',x"3A2A",x"0008");
    gpmc_send('1',x"3A2B",x"0037");
    gpmc_send('1',x"3A2C",x"0007");
    gpmc_send('1',x"3A2D",x"0038");
    gpmc_send('1',x"3A2E",x"0006");
    gpmc_send('1',x"3A2F",x"0039");
    gpmc_send('1',x"3A30",x"0005");
    gpmc_send('1',x"3A31",x"003A");
    gpmc_send('1',x"3A32",x"0004");
    gpmc_send('1',x"3A33",x"003B");
    gpmc_send('1',x"3A34",x"0003");
    gpmc_send('1',x"3A35",x"003C");
    gpmc_send('1',x"3A36",x"0002");
    gpmc_send('1',x"3A37",x"003D");
    gpmc_send('1',x"3A38",x"0001");
    gpmc_send('1',x"3A39",x"003E");
    gpmc_send('1',x"3A3A",x"0000");
    gpmc_send('1',x"3A3B",x"003F");
    gpmc_send('1',x"3A3C",x"0100");
    gpmc_send('1',x"3A3D",x"003E");
    gpmc_send('1',x"3A3E",x"0200");
    gpmc_send('1',x"3A3F",x"003D");
    gpmc_send('1',x"3A40",x"0300");
    gpmc_send('1',x"3A41",x"003C");
    gpmc_send('1',x"3A42",x"0400");
    gpmc_send('1',x"3A43",x"003B");
    gpmc_send('1',x"3A44",x"0500");
    gpmc_send('1',x"3A45",x"003A");
    gpmc_send('1',x"3A46",x"0600");
    gpmc_send('1',x"3A47",x"0039");
    gpmc_send('1',x"3A48",x"0700");
    gpmc_send('1',x"3A49",x"0038");
    gpmc_send('1',x"3A4A",x"0800");
    gpmc_send('1',x"3A4B",x"0037");
    gpmc_send('1',x"3A4C",x"0900");
    gpmc_send('1',x"3A4D",x"0036");
    gpmc_send('1',x"3A4E",x"0A00");
    gpmc_send('1',x"3A4F",x"0035");
    gpmc_send('1',x"3A50",x"0B00");
    gpmc_send('1',x"3A51",x"0034");
    gpmc_send('1',x"3A52",x"0C00");
    gpmc_send('1',x"3A53",x"0033");
    gpmc_send('1',x"3A54",x"0D00");
    gpmc_send('1',x"3A55",x"0032");
    gpmc_send('1',x"3A56",x"0E00");
    gpmc_send('1',x"3A57",x"0031");
    gpmc_send('1',x"3A58",x"0F00");
    gpmc_send('1',x"3A59",x"0030");
    gpmc_send('1',x"3A5A",x"1000");
    gpmc_send('1',x"3A5B",x"002F");
    gpmc_send('1',x"3A5C",x"1100");
    gpmc_send('1',x"3A5D",x"002E");
    gpmc_send('1',x"3A5E",x"1200");
    gpmc_send('1',x"3A5F",x"002D");
    gpmc_send('1',x"3A60",x"1300");
    gpmc_send('1',x"3A61",x"002C");
    gpmc_send('1',x"3A62",x"1400");
    gpmc_send('1',x"3A63",x"002B");
    gpmc_send('1',x"3A64",x"1500");
    gpmc_send('1',x"3A65",x"002A");
    gpmc_send('1',x"3A66",x"1600");
    gpmc_send('1',x"3A67",x"0029");
    gpmc_send('1',x"3A68",x"1700");
    gpmc_send('1',x"3A69",x"0028");
    gpmc_send('1',x"3A6A",x"1800");
    gpmc_send('1',x"3A6B",x"0027");
    gpmc_send('1',x"3A6C",x"1900");
    gpmc_send('1',x"3A6D",x"0026");
    gpmc_send('1',x"3A6E",x"1A00");
    gpmc_send('1',x"3A6F",x"0025");
    gpmc_send('1',x"3A70",x"1B00");
    gpmc_send('1',x"3A71",x"0024");
    gpmc_send('1',x"3A72",x"1C00");
    gpmc_send('1',x"3A73",x"0023");
    gpmc_send('1',x"3A74",x"1D00");
    gpmc_send('1',x"3A75",x"0022");
    gpmc_send('1',x"3A76",x"1E00");
    gpmc_send('1',x"3A77",x"0021");
    gpmc_send('1',x"3A78",x"1F00");
    gpmc_send('1',x"3A79",x"0020");
    gpmc_send('1',x"3A7A",x"2000");
    gpmc_send('1',x"3A7B",x"001F");
    gpmc_send('1',x"3A7C",x"2100");
    gpmc_send('1',x"3A7D",x"001E");
    gpmc_send('1',x"3A7E",x"2200");
    gpmc_send('1',x"3A7F",x"001D");
    gpmc_send('1',x"3A80",x"2300");
    gpmc_send('1',x"3A81",x"001C");
    gpmc_send('1',x"3A82",x"2400");
    gpmc_send('1',x"3A83",x"001B");
    gpmc_send('1',x"3A84",x"2500");
    gpmc_send('1',x"3A85",x"001A");
    gpmc_send('1',x"3A86",x"2600");
    gpmc_send('1',x"3A87",x"0019");
    gpmc_send('1',x"3A88",x"2700");
    gpmc_send('1',x"3A89",x"0018");
    gpmc_send('1',x"3A8A",x"2800");
    gpmc_send('1',x"3A8B",x"0017");
    gpmc_send('1',x"3A8C",x"2900");
    gpmc_send('1',x"3A8D",x"0016");
    gpmc_send('1',x"3A8E",x"2A00");
    gpmc_send('1',x"3A8F",x"0015");
    gpmc_send('1',x"3A90",x"2B00");
    gpmc_send('1',x"3A91",x"0014");
    gpmc_send('1',x"3A92",x"2C00");
    gpmc_send('1',x"3A93",x"0013");
    gpmc_send('1',x"3A94",x"2D00");
    gpmc_send('1',x"3A95",x"0012");
    gpmc_send('1',x"3A96",x"2E00");
    gpmc_send('1',x"3A97",x"0011");
    gpmc_send('1',x"3A98",x"2F00");
    gpmc_send('1',x"3A99",x"0010");
    gpmc_send('1',x"3A9A",x"3000");
    gpmc_send('1',x"3A9B",x"000F");
    gpmc_send('1',x"3A9C",x"3100");
    gpmc_send('1',x"3A9D",x"000E");
    gpmc_send('1',x"3A9E",x"3200");
    gpmc_send('1',x"3A9F",x"000D");
    gpmc_send('1',x"3AA0",x"3300");
    gpmc_send('1',x"3AA1",x"000C");
    gpmc_send('1',x"3AA2",x"3400");
    gpmc_send('1',x"3AA3",x"000B");
    gpmc_send('1',x"3AA4",x"3500");
    gpmc_send('1',x"3AA5",x"000A");
    gpmc_send('1',x"3AA6",x"3600");
    gpmc_send('1',x"3AA7",x"0009");
    gpmc_send('1',x"3AA8",x"3700");
    gpmc_send('1',x"3AA9",x"0008");
    gpmc_send('1',x"3AAA",x"3800");
    gpmc_send('1',x"3AAB",x"0007");
    gpmc_send('1',x"3AAC",x"3900");
    gpmc_send('1',x"3AAD",x"0006");
    gpmc_send('1',x"3AAE",x"3A00");
    gpmc_send('1',x"3AAF",x"0005");
    gpmc_send('1',x"3AB0",x"3B00");
    gpmc_send('1',x"3AB1",x"0004");
    gpmc_send('1',x"3AB2",x"3C00");
    gpmc_send('1',x"3AB3",x"0003");
    gpmc_send('1',x"3AB4",x"3D00");
    gpmc_send('1',x"3AB5",x"0002");
    gpmc_send('1',x"3AB6",x"3E00");
    gpmc_send('1',x"3AB7",x"0001");
    gpmc_send('1',x"3AB8",x"3F00");
    gpmc_send('1',x"3AB9",x"0000");
    gpmc_send('1',x"3ABA",x"3F01");
    gpmc_send('1',x"3ABB",x"0000");
    gpmc_send('1',x"3ABC",x"3E02");
    gpmc_send('1',x"3ABD",x"0000");
    gpmc_send('1',x"3ABE",x"3D03");
    gpmc_send('1',x"3ABF",x"0000");
    gpmc_send('1',x"3AC0",x"3C04");
    gpmc_send('1',x"3AC1",x"0000");
    gpmc_send('1',x"3AC2",x"3B05");
    gpmc_send('1',x"3AC3",x"0000");
    gpmc_send('1',x"3AC4",x"3A06");
    gpmc_send('1',x"3AC5",x"0000");
    gpmc_send('1',x"3AC6",x"3907");
    gpmc_send('1',x"3AC7",x"0000");
    gpmc_send('1',x"3AC8",x"3808");
    gpmc_send('1',x"3AC9",x"0000");
    gpmc_send('1',x"3ACA",x"3709");
    gpmc_send('1',x"3ACB",x"0000");
    gpmc_send('1',x"3ACC",x"360A");
    gpmc_send('1',x"3ACD",x"0000");
    gpmc_send('1',x"3ACE",x"350B");
    gpmc_send('1',x"3ACF",x"0000");
    gpmc_send('1',x"3AD0",x"340C");
    gpmc_send('1',x"3AD1",x"0000");
    gpmc_send('1',x"3AD2",x"330D");
    gpmc_send('1',x"3AD3",x"0000");
    gpmc_send('1',x"3AD4",x"320E");
    gpmc_send('1',x"3AD5",x"0000");
    gpmc_send('1',x"3AD6",x"310F");
    gpmc_send('1',x"3AD7",x"0000");
    gpmc_send('1',x"3AD8",x"3010");
    gpmc_send('1',x"3AD9",x"0000");
    gpmc_send('1',x"3ADA",x"2F11");
    gpmc_send('1',x"3ADB",x"0000");
    gpmc_send('1',x"3ADC",x"2E12");
    gpmc_send('1',x"3ADD",x"0000");
    gpmc_send('1',x"3ADE",x"2D13");
    gpmc_send('1',x"3ADF",x"0000");
    gpmc_send('1',x"3AE0",x"2C14");
    gpmc_send('1',x"3AE1",x"0000");
    gpmc_send('1',x"3AE2",x"2B15");
    gpmc_send('1',x"3AE3",x"0000");
    gpmc_send('1',x"3AE4",x"2A16");
    gpmc_send('1',x"3AE5",x"0000");
    gpmc_send('1',x"3AE6",x"2917");
    gpmc_send('1',x"3AE7",x"0000");
    gpmc_send('1',x"3AE8",x"2818");
    gpmc_send('1',x"3AE9",x"0000");
    gpmc_send('1',x"3AEA",x"2719");
    gpmc_send('1',x"3AEB",x"0000");
    gpmc_send('1',x"3AEC",x"261A");
    gpmc_send('1',x"3AED",x"0000");
    gpmc_send('1',x"3AEE",x"251B");
    gpmc_send('1',x"3AEF",x"0000");
    gpmc_send('1',x"3AF0",x"241C");
    gpmc_send('1',x"3AF1",x"0000");
    gpmc_send('1',x"3AF2",x"231D");
    gpmc_send('1',x"3AF3",x"0000");
    gpmc_send('1',x"3AF4",x"221E");
    gpmc_send('1',x"3AF5",x"0000");
    gpmc_send('1',x"3AF6",x"211F");
    gpmc_send('1',x"3AF7",x"0000");
    gpmc_send('1',x"3AF8",x"2020");
    gpmc_send('1',x"3AF9",x"0000");
    gpmc_send('1',x"3AFA",x"1F21");
    gpmc_send('1',x"3AFB",x"0000");
    gpmc_send('1',x"3AFC",x"1E22");
    gpmc_send('1',x"3AFD",x"0000");
    gpmc_send('1',x"3AFE",x"1D23");
    gpmc_send('1',x"3AFF",x"0000");
    gpmc_send('1',x"3B00",x"1C24");
    gpmc_send('1',x"3B01",x"0000");
    gpmc_send('1',x"3B02",x"1B25");
    gpmc_send('1',x"3B03",x"0000");
    gpmc_send('1',x"3B04",x"1A26");
    gpmc_send('1',x"3B05",x"0000");
    gpmc_send('1',x"3B06",x"1927");
    gpmc_send('1',x"3B07",x"0000");
    gpmc_send('1',x"3B08",x"1828");
    gpmc_send('1',x"3B09",x"0000");
    gpmc_send('1',x"3B0A",x"1729");
    gpmc_send('1',x"3B0B",x"0000");
    gpmc_send('1',x"3B0C",x"162A");
    gpmc_send('1',x"3B0D",x"0000");
    gpmc_send('1',x"3B0E",x"152B");
    gpmc_send('1',x"3B0F",x"0000");
    gpmc_send('1',x"3B10",x"142C");
    gpmc_send('1',x"3B11",x"0000");
    gpmc_send('1',x"3B12",x"132D");
    gpmc_send('1',x"3B13",x"0000");
    gpmc_send('1',x"3B14",x"122E");
    gpmc_send('1',x"3B15",x"0000");
    gpmc_send('1',x"3B16",x"112F");
    gpmc_send('1',x"3B17",x"0000");
    gpmc_send('1',x"3B18",x"1030");
    gpmc_send('1',x"3B19",x"0000");
    gpmc_send('1',x"3B1A",x"0F31");
    gpmc_send('1',x"3B1B",x"0000");
    gpmc_send('1',x"3B1C",x"0E32");
    gpmc_send('1',x"3B1D",x"0000");
    gpmc_send('1',x"3B1E",x"0D33");
    gpmc_send('1',x"3B1F",x"0000");
    gpmc_send('1',x"3B20",x"0C34");
    gpmc_send('1',x"3B21",x"0000");
    gpmc_send('1',x"3B22",x"0B35");
    gpmc_send('1',x"3B23",x"0000");
    gpmc_send('1',x"3B24",x"0A36");
    gpmc_send('1',x"3B25",x"0000");
    gpmc_send('1',x"3B26",x"0937");
    gpmc_send('1',x"3B27",x"0000");
    gpmc_send('1',x"3B28",x"0838");
    gpmc_send('1',x"3B29",x"0000");
    gpmc_send('1',x"3B2A",x"0739");
    gpmc_send('1',x"3B2B",x"0000");
    gpmc_send('1',x"3B2C",x"063A");
    gpmc_send('1',x"3B2D",x"0000");
    gpmc_send('1',x"3B2E",x"053B");
    gpmc_send('1',x"3B2F",x"0000");
    gpmc_send('1',x"3B30",x"043C");
    gpmc_send('1',x"3B31",x"0000");
    gpmc_send('1',x"3B32",x"033D");
    gpmc_send('1',x"3B33",x"0000");
    gpmc_send('1',x"3B34",x"023E");
    gpmc_send('1',x"3B35",x"0000");
    gpmc_send('1',x"3B36",x"013F");
    gpmc_send('1',x"3B37",x"0000");
    gpmc_send('1',x"3B38",x"003F");
    gpmc_send('1',x"3B39",x"0000");
    gpmc_send('1',x"3B3A",x"003E");
    gpmc_send('1',x"3B3B",x"0001");
    gpmc_send('1',x"3B3C",x"003D");
    gpmc_send('1',x"3B3D",x"0002");
    gpmc_send('1',x"3B3E",x"003C");
    gpmc_send('1',x"3B3F",x"0003");
    gpmc_send('1',x"3B40",x"003B");
    gpmc_send('1',x"3B41",x"0004");
    gpmc_send('1',x"3B42",x"003A");
    gpmc_send('1',x"3B43",x"0005");
    gpmc_send('1',x"3B44",x"0039");
    gpmc_send('1',x"3B45",x"0006");
    gpmc_send('1',x"3B46",x"0038");
    gpmc_send('1',x"3B47",x"0007");
    gpmc_send('1',x"3B48",x"0037");
    gpmc_send('1',x"3B49",x"0008");
    gpmc_send('1',x"3B4A",x"0036");
    gpmc_send('1',x"3B4B",x"0009");
    gpmc_send('1',x"3B4C",x"0035");
    gpmc_send('1',x"3B4D",x"000A");
    gpmc_send('1',x"3B4E",x"0034");
    gpmc_send('1',x"3B4F",x"000B");
    gpmc_send('1',x"3B50",x"0033");
    gpmc_send('1',x"3B51",x"000C");
    gpmc_send('1',x"3B52",x"0032");
    gpmc_send('1',x"3B53",x"000D");
    gpmc_send('1',x"3B54",x"0031");
    gpmc_send('1',x"3B55",x"000E");
    gpmc_send('1',x"3B56",x"0030");
    gpmc_send('1',x"3B57",x"000F");
    gpmc_send('1',x"3B58",x"002F");
    gpmc_send('1',x"3B59",x"0010");
    gpmc_send('1',x"3B5A",x"002E");
    gpmc_send('1',x"3B5B",x"0011");
    gpmc_send('1',x"3B5C",x"002D");
    gpmc_send('1',x"3B5D",x"0012");
    gpmc_send('1',x"3B5E",x"002C");
    gpmc_send('1',x"3B5F",x"0013");
    gpmc_send('1',x"3B60",x"002B");
    gpmc_send('1',x"3B61",x"0014");
    gpmc_send('1',x"3B62",x"002A");
    gpmc_send('1',x"3B63",x"0015");
    gpmc_send('1',x"3B64",x"0029");
    gpmc_send('1',x"3B65",x"0016");
    gpmc_send('1',x"3B66",x"0028");
    gpmc_send('1',x"3B67",x"0017");
    gpmc_send('1',x"3B68",x"0027");
    gpmc_send('1',x"3B69",x"0018");
    gpmc_send('1',x"3B6A",x"0026");
    gpmc_send('1',x"3B6B",x"0019");
    gpmc_send('1',x"3B6C",x"0025");
    gpmc_send('1',x"3B6D",x"001A");
    gpmc_send('1',x"3B6E",x"0024");
    gpmc_send('1',x"3B6F",x"001B");
    gpmc_send('1',x"3B70",x"0023");
    gpmc_send('1',x"3B71",x"001C");
    gpmc_send('1',x"3B72",x"0022");
    gpmc_send('1',x"3B73",x"001D");
    gpmc_send('1',x"3B74",x"0021");
    gpmc_send('1',x"3B75",x"001E");
    gpmc_send('1',x"3B76",x"0020");
    gpmc_send('1',x"3B77",x"001F");
    gpmc_send('1',x"3B78",x"001F");
    gpmc_send('1',x"3B79",x"0020");
    gpmc_send('1',x"3B7A",x"001E");
    gpmc_send('1',x"3B7B",x"0021");
    gpmc_send('1',x"3B7C",x"001D");
    gpmc_send('1',x"3B7D",x"0022");
    gpmc_send('1',x"3B7E",x"001C");
    gpmc_send('1',x"3B7F",x"0023");
    gpmc_send('1',x"3B80",x"001B");
    gpmc_send('1',x"3B81",x"0024");
    gpmc_send('1',x"3B82",x"001A");
    gpmc_send('1',x"3B83",x"0025");
    gpmc_send('1',x"3B84",x"0019");
    gpmc_send('1',x"3B85",x"0026");
    gpmc_send('1',x"3B86",x"0018");
    gpmc_send('1',x"3B87",x"0027");
    gpmc_send('1',x"3B88",x"0017");
    gpmc_send('1',x"3B89",x"0028");
    gpmc_send('1',x"3B8A",x"0016");
    gpmc_send('1',x"3B8B",x"0029");
    gpmc_send('1',x"3B8C",x"0015");
    gpmc_send('1',x"3B8D",x"002A");
    gpmc_send('1',x"3B8E",x"0014");
    gpmc_send('1',x"3B8F",x"002B");
    gpmc_send('1',x"3B90",x"0013");
    gpmc_send('1',x"3B91",x"002C");
    gpmc_send('1',x"3B92",x"0012");
    gpmc_send('1',x"3B93",x"002D");
    gpmc_send('1',x"3B94",x"0011");
    gpmc_send('1',x"3B95",x"002E");
    gpmc_send('1',x"3B96",x"0010");
    gpmc_send('1',x"3B97",x"002F");
    gpmc_send('1',x"3B98",x"000F");
    gpmc_send('1',x"3B99",x"0030");
    gpmc_send('1',x"3B9A",x"000E");
    gpmc_send('1',x"3B9B",x"0031");
    gpmc_send('1',x"3B9C",x"000D");
    gpmc_send('1',x"3B9D",x"0032");
    gpmc_send('1',x"3B9E",x"000C");
    gpmc_send('1',x"3B9F",x"0033");
    gpmc_send('1',x"3BA0",x"000B");
    gpmc_send('1',x"3BA1",x"0034");
    gpmc_send('1',x"3BA2",x"000A");
    gpmc_send('1',x"3BA3",x"0035");
    gpmc_send('1',x"3BA4",x"0009");
    gpmc_send('1',x"3BA5",x"0036");
    gpmc_send('1',x"3BA6",x"0008");
    gpmc_send('1',x"3BA7",x"0037");
    gpmc_send('1',x"3BA8",x"0007");
    gpmc_send('1',x"3BA9",x"0038");
    gpmc_send('1',x"3BAA",x"0006");
    gpmc_send('1',x"3BAB",x"0039");
    gpmc_send('1',x"3BAC",x"0005");
    gpmc_send('1',x"3BAD",x"003A");
    gpmc_send('1',x"3BAE",x"0004");
    gpmc_send('1',x"3BAF",x"003B");
    gpmc_send('1',x"3BB0",x"0003");
    gpmc_send('1',x"3BB1",x"003C");
    gpmc_send('1',x"3BB2",x"0002");
    gpmc_send('1',x"3BB3",x"003D");
    gpmc_send('1',x"3BB4",x"0001");
    gpmc_send('1',x"3BB5",x"003E");
    gpmc_send('1',x"3BB6",x"0000");
    gpmc_send('1',x"3BB7",x"003F");
    gpmc_send('1',x"3BB8",x"0100");
    gpmc_send('1',x"3BB9",x"003E");
    gpmc_send('1',x"3BBA",x"0200");
    gpmc_send('1',x"3BBB",x"003D");
    gpmc_send('1',x"3BBC",x"0300");
    gpmc_send('1',x"3BBD",x"003C");
    gpmc_send('1',x"3BBE",x"0400");
    gpmc_send('1',x"3BBF",x"003B");
    gpmc_send('1',x"3BC0",x"0500");
    gpmc_send('1',x"3BC1",x"003A");
    gpmc_send('1',x"3BC2",x"0600");
    gpmc_send('1',x"3BC3",x"0039");
    gpmc_send('1',x"3BC4",x"0700");
    gpmc_send('1',x"3BC5",x"0038");
    gpmc_send('1',x"3BC6",x"0800");
    gpmc_send('1',x"3BC7",x"0037");
    gpmc_send('1',x"3BC8",x"0900");
    gpmc_send('1',x"3BC9",x"0036");
    gpmc_send('1',x"3BCA",x"0A00");
    gpmc_send('1',x"3BCB",x"0035");
    gpmc_send('1',x"3BCC",x"0B00");
    gpmc_send('1',x"3BCD",x"0034");
    gpmc_send('1',x"3BCE",x"0C00");
    gpmc_send('1',x"3BCF",x"0033");
    gpmc_send('1',x"3BD0",x"0D00");
    gpmc_send('1',x"3BD1",x"0032");
    gpmc_send('1',x"3BD2",x"0E00");
    gpmc_send('1',x"3BD3",x"0031");
    gpmc_send('1',x"3BD4",x"0F00");
    gpmc_send('1',x"3BD5",x"0030");
    gpmc_send('1',x"3BD6",x"1000");
    gpmc_send('1',x"3BD7",x"002F");
    gpmc_send('1',x"3BD8",x"1100");
    gpmc_send('1',x"3BD9",x"002E");
    gpmc_send('1',x"3BDA",x"1200");
    gpmc_send('1',x"3BDB",x"002D");
    gpmc_send('1',x"3BDC",x"1300");
    gpmc_send('1',x"3BDD",x"002C");
    gpmc_send('1',x"3BDE",x"1400");
    gpmc_send('1',x"3BDF",x"002B");
    gpmc_send('1',x"3BE0",x"1500");
    gpmc_send('1',x"3BE1",x"002A");
    gpmc_send('1',x"3BE2",x"1600");
    gpmc_send('1',x"3BE3",x"0029");
    gpmc_send('1',x"3BE4",x"1700");
    gpmc_send('1',x"3BE5",x"0028");
    gpmc_send('1',x"3BE6",x"1800");
    gpmc_send('1',x"3BE7",x"0027");
    gpmc_send('1',x"3BE8",x"1900");
    gpmc_send('1',x"3BE9",x"0026");
    gpmc_send('1',x"3BEA",x"1A00");
    gpmc_send('1',x"3BEB",x"0025");
    gpmc_send('1',x"3BEC",x"1B00");
    gpmc_send('1',x"3BED",x"0024");
    gpmc_send('1',x"3BEE",x"1C00");
    gpmc_send('1',x"3BEF",x"0023");
    gpmc_send('1',x"3BF0",x"1D00");
    gpmc_send('1',x"3BF1",x"0022");
    gpmc_send('1',x"3BF2",x"1E00");
    gpmc_send('1',x"3BF3",x"0021");
    gpmc_send('1',x"3BF4",x"1F00");
    gpmc_send('1',x"3BF5",x"0020");
    gpmc_send('1',x"3BF6",x"2000");
    gpmc_send('1',x"3BF7",x"001F");
    gpmc_send('1',x"3BF8",x"2100");
    gpmc_send('1',x"3BF9",x"001E");
    gpmc_send('1',x"3BFA",x"2200");
    gpmc_send('1',x"3BFB",x"001D");
    gpmc_send('1',x"3BFC",x"2300");
    gpmc_send('1',x"3BFD",x"001C");
    gpmc_send('1',x"3BFE",x"2400");
    gpmc_send('1',x"3BFF",x"001B");
    gpmc_send('1',x"3C00",x"2500");
    gpmc_send('1',x"3C01",x"001A");
    gpmc_send('1',x"3C02",x"2600");
    gpmc_send('1',x"3C03",x"0019");
    gpmc_send('1',x"3C04",x"2700");
    gpmc_send('1',x"3C05",x"0018");
    gpmc_send('1',x"3C06",x"2800");
    gpmc_send('1',x"3C07",x"0017");
    gpmc_send('1',x"3C08",x"2900");
    gpmc_send('1',x"3C09",x"0016");
    gpmc_send('1',x"3C0A",x"2A00");
    gpmc_send('1',x"3C0B",x"0015");
    gpmc_send('1',x"3C0C",x"2B00");
    gpmc_send('1',x"3C0D",x"0014");
    gpmc_send('1',x"3C0E",x"2C00");
    gpmc_send('1',x"3C0F",x"0013");
    gpmc_send('1',x"3C10",x"2D00");
    gpmc_send('1',x"3C11",x"0012");
    gpmc_send('1',x"3C12",x"2E00");
    gpmc_send('1',x"3C13",x"0011");
    gpmc_send('1',x"3C14",x"2F00");
    gpmc_send('1',x"3C15",x"0010");
    gpmc_send('1',x"3C16",x"3000");
    gpmc_send('1',x"3C17",x"000F");
    gpmc_send('1',x"3C18",x"3100");
    gpmc_send('1',x"3C19",x"000E");
    gpmc_send('1',x"3C1A",x"3200");
    gpmc_send('1',x"3C1B",x"000D");
    gpmc_send('1',x"3C1C",x"3300");
    gpmc_send('1',x"3C1D",x"000C");
    gpmc_send('1',x"3C1E",x"3400");
    gpmc_send('1',x"3C1F",x"000B");
    gpmc_send('1',x"3C20",x"3500");
    gpmc_send('1',x"3C21",x"000A");
    gpmc_send('1',x"3C22",x"3600");
    gpmc_send('1',x"3C23",x"0009");
    gpmc_send('1',x"3C24",x"3700");
    gpmc_send('1',x"3C25",x"0008");
    gpmc_send('1',x"3C26",x"3800");
    gpmc_send('1',x"3C27",x"0007");
    gpmc_send('1',x"3C28",x"3900");
    gpmc_send('1',x"3C29",x"0006");
    gpmc_send('1',x"3C2A",x"3A00");
    gpmc_send('1',x"3C2B",x"0005");
    gpmc_send('1',x"3C2C",x"3B00");
    gpmc_send('1',x"3C2D",x"0004");
    gpmc_send('1',x"3C2E",x"3C00");
    gpmc_send('1',x"3C2F",x"0003");
    gpmc_send('1',x"3C30",x"3D00");
    gpmc_send('1',x"3C31",x"0002");
    gpmc_send('1',x"3C32",x"3E00");
    gpmc_send('1',x"3C33",x"0001");
    gpmc_send('1',x"3C34",x"3F00");
    gpmc_send('1',x"3C35",x"0000");
    gpmc_send('1',x"3C36",x"3F01");
    gpmc_send('1',x"3C37",x"0000");
    gpmc_send('1',x"3C38",x"3E02");
    gpmc_send('1',x"3C39",x"0000");
    gpmc_send('1',x"3C3A",x"3D03");
    gpmc_send('1',x"3C3B",x"0000");
    gpmc_send('1',x"3C3C",x"3C04");
    gpmc_send('1',x"3C3D",x"0000");
    gpmc_send('1',x"3C3E",x"3B05");
    gpmc_send('1',x"3C3F",x"0000");
    gpmc_send('1',x"3C40",x"3A06");
    gpmc_send('1',x"3C41",x"0000");
    gpmc_send('1',x"3C42",x"3907");
    gpmc_send('1',x"3C43",x"0000");
    gpmc_send('1',x"3C44",x"3808");
    gpmc_send('1',x"3C45",x"0000");
    gpmc_send('1',x"3C46",x"3709");
    gpmc_send('1',x"3C47",x"0000");
    gpmc_send('1',x"3C48",x"360A");
    gpmc_send('1',x"3C49",x"0000");
    gpmc_send('1',x"3C4A",x"350B");
    gpmc_send('1',x"3C4B",x"0000");
    gpmc_send('1',x"3C4C",x"340C");
    gpmc_send('1',x"3C4D",x"0000");
    gpmc_send('1',x"3C4E",x"330D");
    gpmc_send('1',x"3C4F",x"0000");
    gpmc_send('1',x"3C50",x"320E");
    gpmc_send('1',x"3C51",x"0000");
    gpmc_send('1',x"3C52",x"310F");
    gpmc_send('1',x"3C53",x"0000");
    gpmc_send('1',x"3C54",x"3010");
    gpmc_send('1',x"3C55",x"0000");
    gpmc_send('1',x"3C56",x"2F11");
    gpmc_send('1',x"3C57",x"0000");
    gpmc_send('1',x"3C58",x"2E12");
    gpmc_send('1',x"3C59",x"0000");
    gpmc_send('1',x"3C5A",x"2D13");
    gpmc_send('1',x"3C5B",x"0000");
    gpmc_send('1',x"3C5C",x"2C14");
    gpmc_send('1',x"3C5D",x"0000");
    gpmc_send('1',x"3C5E",x"2B15");
    gpmc_send('1',x"3C5F",x"0000");
    gpmc_send('1',x"3C60",x"2A16");
    gpmc_send('1',x"3C61",x"0000");
    gpmc_send('1',x"3C62",x"2917");
    gpmc_send('1',x"3C63",x"0000");
    gpmc_send('1',x"3C64",x"2818");
    gpmc_send('1',x"3C65",x"0000");
    gpmc_send('1',x"3C66",x"2719");
    gpmc_send('1',x"3C67",x"0000");
    gpmc_send('1',x"3C68",x"261A");
    gpmc_send('1',x"3C69",x"0000");
    gpmc_send('1',x"3C6A",x"251B");
    gpmc_send('1',x"3C6B",x"0000");
    gpmc_send('1',x"3C6C",x"241C");
    gpmc_send('1',x"3C6D",x"0000");
    gpmc_send('1',x"3C6E",x"231D");
    gpmc_send('1',x"3C6F",x"0000");
    gpmc_send('1',x"3C70",x"221E");
    gpmc_send('1',x"3C71",x"0000");
    gpmc_send('1',x"3C72",x"211F");
    gpmc_send('1',x"3C73",x"0000");
    gpmc_send('1',x"3C74",x"2020");
    gpmc_send('1',x"3C75",x"0000");
    gpmc_send('1',x"3C76",x"1F21");
    gpmc_send('1',x"3C77",x"0000");
    gpmc_send('1',x"3C78",x"1E22");
    gpmc_send('1',x"3C79",x"0000");
    gpmc_send('1',x"3C7A",x"1D23");
    gpmc_send('1',x"3C7B",x"0000");
    gpmc_send('1',x"3C7C",x"1C24");
    gpmc_send('1',x"3C7D",x"0000");
    gpmc_send('1',x"3C7E",x"1B25");
    gpmc_send('1',x"3C7F",x"0000");
    gpmc_send('1',x"3C80",x"1A26");
    gpmc_send('1',x"3C81",x"0000");
    gpmc_send('1',x"3C82",x"1927");
    gpmc_send('1',x"3C83",x"0000");
    gpmc_send('1',x"3C84",x"1828");
    gpmc_send('1',x"3C85",x"0000");
    gpmc_send('1',x"3C86",x"1729");
    gpmc_send('1',x"3C87",x"0000");
    gpmc_send('1',x"3C88",x"162A");
    gpmc_send('1',x"3C89",x"0000");
    gpmc_send('1',x"3C8A",x"152B");
    gpmc_send('1',x"3C8B",x"0000");
    gpmc_send('1',x"3C8C",x"142C");
    gpmc_send('1',x"3C8D",x"0000");
    gpmc_send('1',x"3C8E",x"132D");
    gpmc_send('1',x"3C8F",x"0000");
    gpmc_send('1',x"3C90",x"122E");
    gpmc_send('1',x"3C91",x"0000");
    gpmc_send('1',x"3C92",x"112F");
    gpmc_send('1',x"3C93",x"0000");
    gpmc_send('1',x"3C94",x"1030");
    gpmc_send('1',x"3C95",x"0000");
    gpmc_send('1',x"3C96",x"0F31");
    gpmc_send('1',x"3C97",x"0000");
    gpmc_send('1',x"3C98",x"0E32");
    gpmc_send('1',x"3C99",x"0000");
    gpmc_send('1',x"3C9A",x"0D33");
    gpmc_send('1',x"3C9B",x"0000");
    gpmc_send('1',x"3C9C",x"0C34");
    gpmc_send('1',x"3C9D",x"0000");
    gpmc_send('1',x"3C9E",x"0B35");
    gpmc_send('1',x"3C9F",x"0000");
    gpmc_send('1',x"3CA0",x"0A36");
    gpmc_send('1',x"3CA1",x"0000");
    gpmc_send('1',x"3CA2",x"0937");
    gpmc_send('1',x"3CA3",x"0000");
    gpmc_send('1',x"3CA4",x"0838");
    gpmc_send('1',x"3CA5",x"0000");
    gpmc_send('1',x"3CA6",x"0739");
    gpmc_send('1',x"3CA7",x"0000");
    gpmc_send('1',x"3CA8",x"063A");
    gpmc_send('1',x"3CA9",x"0000");
    gpmc_send('1',x"3CAA",x"053B");
    gpmc_send('1',x"3CAB",x"0000");
    gpmc_send('1',x"3CAC",x"043C");
    gpmc_send('1',x"3CAD",x"0000");
    gpmc_send('1',x"3CAE",x"033D");
    gpmc_send('1',x"3CAF",x"0000");
    gpmc_send('1',x"3CB0",x"023E");
    gpmc_send('1',x"3CB1",x"0000");
    gpmc_send('1',x"3CB2",x"013F");
    gpmc_send('1',x"3CB3",x"0000");
    gpmc_send('1',x"3CB4",x"003F");
    gpmc_send('1',x"3CB5",x"0000");
    gpmc_send('1',x"3CB6",x"003E");
    gpmc_send('1',x"3CB7",x"0001");
    gpmc_send('1',x"3CB8",x"003D");
    gpmc_send('1',x"3CB9",x"0002");
    gpmc_send('1',x"3CBA",x"003C");
    gpmc_send('1',x"3CBB",x"0003");
    gpmc_send('1',x"3CBC",x"003B");
    gpmc_send('1',x"3CBD",x"0004");
    gpmc_send('1',x"3CBE",x"003A");
    gpmc_send('1',x"3CBF",x"0005");
    gpmc_send('1',x"3CC0",x"0039");
    gpmc_send('1',x"3CC1",x"0006");
    gpmc_send('1',x"3CC2",x"0038");
    gpmc_send('1',x"3CC3",x"0007");
    gpmc_send('1',x"3CC4",x"0037");
    gpmc_send('1',x"3CC5",x"0008");
    gpmc_send('1',x"3CC6",x"0036");
    gpmc_send('1',x"3CC7",x"0009");
    gpmc_send('1',x"3CC8",x"0035");
    gpmc_send('1',x"3CC9",x"000A");
    gpmc_send('1',x"3CCA",x"0034");
    gpmc_send('1',x"3CCB",x"000B");
    gpmc_send('1',x"3CCC",x"0033");
    gpmc_send('1',x"3CCD",x"000C");
    gpmc_send('1',x"3CCE",x"0032");
    gpmc_send('1',x"3CCF",x"000D");
    gpmc_send('1',x"3CD0",x"0031");
    gpmc_send('1',x"3CD1",x"000E");
    gpmc_send('1',x"3CD2",x"0030");
    gpmc_send('1',x"3CD3",x"000F");
    gpmc_send('1',x"3CD4",x"002F");
    gpmc_send('1',x"3CD5",x"0010");
    gpmc_send('1',x"3CD6",x"002E");
    gpmc_send('1',x"3CD7",x"0011");
    gpmc_send('1',x"3CD8",x"002D");
    gpmc_send('1',x"3CD9",x"0012");
    gpmc_send('1',x"3CDA",x"002C");
    gpmc_send('1',x"3CDB",x"0013");
    gpmc_send('1',x"3CDC",x"002B");
    gpmc_send('1',x"3CDD",x"0014");
    gpmc_send('1',x"3CDE",x"002A");
    gpmc_send('1',x"3CDF",x"0015");
    gpmc_send('1',x"3CE0",x"0029");
    gpmc_send('1',x"3CE1",x"0016");
    gpmc_send('1',x"3CE2",x"0028");
    gpmc_send('1',x"3CE3",x"0017");
    gpmc_send('1',x"3CE4",x"0027");
    gpmc_send('1',x"3CE5",x"0018");
    gpmc_send('1',x"3CE6",x"0026");
    gpmc_send('1',x"3CE7",x"0019");
    gpmc_send('1',x"3CE8",x"0025");
    gpmc_send('1',x"3CE9",x"001A");
    gpmc_send('1',x"3CEA",x"0024");
    gpmc_send('1',x"3CEB",x"001B");
    gpmc_send('1',x"3CEC",x"0023");
    gpmc_send('1',x"3CED",x"001C");
    gpmc_send('1',x"3CEE",x"0022");
    gpmc_send('1',x"3CEF",x"001D");
    gpmc_send('1',x"3CF0",x"0021");
    gpmc_send('1',x"3CF1",x"001E");
    gpmc_send('1',x"3CF2",x"0020");
    gpmc_send('1',x"3CF3",x"001F");
    gpmc_send('1',x"3CF4",x"001F");
    gpmc_send('1',x"3CF5",x"0020");
    gpmc_send('1',x"3CF6",x"001E");
    gpmc_send('1',x"3CF7",x"0021");
    gpmc_send('1',x"3CF8",x"001D");
    gpmc_send('1',x"3CF9",x"0022");
    gpmc_send('1',x"3CFA",x"001C");
    gpmc_send('1',x"3CFB",x"0023");
    gpmc_send('1',x"3CFC",x"001B");
    gpmc_send('1',x"3CFD",x"0024");
    gpmc_send('1',x"3CFE",x"001A");
    gpmc_send('1',x"3CFF",x"0025");
    gpmc_send('1',x"3D00",x"0019");
    gpmc_send('1',x"3D01",x"0026");
    gpmc_send('1',x"3D02",x"0018");
    gpmc_send('1',x"3D03",x"0027");
    gpmc_send('1',x"3D04",x"0017");
    gpmc_send('1',x"3D05",x"0028");
    gpmc_send('1',x"3D06",x"0016");
    gpmc_send('1',x"3D07",x"0029");
    gpmc_send('1',x"3D08",x"0015");
    gpmc_send('1',x"3D09",x"002A");
    gpmc_send('1',x"3D0A",x"0014");
    gpmc_send('1',x"3D0B",x"002B");
    gpmc_send('1',x"3D0C",x"0013");
    gpmc_send('1',x"3D0D",x"002C");
    gpmc_send('1',x"3D0E",x"0012");
    gpmc_send('1',x"3D0F",x"002D");
    gpmc_send('1',x"3D10",x"0011");
    gpmc_send('1',x"3D11",x"002E");
    gpmc_send('1',x"3D12",x"0010");
    gpmc_send('1',x"3D13",x"002F");
    gpmc_send('1',x"3D14",x"000F");
    gpmc_send('1',x"3D15",x"0030");
    gpmc_send('1',x"3D16",x"000E");
    gpmc_send('1',x"3D17",x"0031");
    gpmc_send('1',x"3D18",x"000D");
    gpmc_send('1',x"3D19",x"0032");
    gpmc_send('1',x"3D1A",x"000C");
    gpmc_send('1',x"3D1B",x"0033");
    gpmc_send('1',x"3D1C",x"000B");
    gpmc_send('1',x"3D1D",x"0034");
    gpmc_send('1',x"3D1E",x"000A");
    gpmc_send('1',x"3D1F",x"0035");
    gpmc_send('1',x"3D20",x"0009");
    gpmc_send('1',x"3D21",x"0036");
    gpmc_send('1',x"3D22",x"0008");
    gpmc_send('1',x"3D23",x"0037");
    gpmc_send('1',x"3D24",x"0007");
    gpmc_send('1',x"3D25",x"0038");
    gpmc_send('1',x"3D26",x"0006");
    gpmc_send('1',x"3D27",x"0039");
    gpmc_send('1',x"3D28",x"0005");
    gpmc_send('1',x"3D29",x"003A");
    gpmc_send('1',x"3D2A",x"0004");
    gpmc_send('1',x"3D2B",x"003B");
    gpmc_send('1',x"3D2C",x"0003");
    gpmc_send('1',x"3D2D",x"003C");
    gpmc_send('1',x"3D2E",x"0002");
    gpmc_send('1',x"3D2F",x"003D");
    gpmc_send('1',x"3D30",x"0001");
    gpmc_send('1',x"3D31",x"003E");
    gpmc_send('1',x"3D32",x"0000");
    gpmc_send('1',x"3D33",x"003F");
    gpmc_send('1',x"3D34",x"0100");
    gpmc_send('1',x"3D35",x"003E");
    gpmc_send('1',x"3D36",x"0200");
    gpmc_send('1',x"3D37",x"003D");
    gpmc_send('1',x"3D38",x"0300");
    gpmc_send('1',x"3D39",x"003C");
    gpmc_send('1',x"3D3A",x"0400");
    gpmc_send('1',x"3D3B",x"003B");
    gpmc_send('1',x"3D3C",x"0500");
    gpmc_send('1',x"3D3D",x"003A");
    gpmc_send('1',x"3D3E",x"0600");
    gpmc_send('1',x"3D3F",x"0039");
    gpmc_send('1',x"3D40",x"0700");
    gpmc_send('1',x"3D41",x"0038");
    gpmc_send('1',x"3D42",x"0800");
    gpmc_send('1',x"3D43",x"0037");
    gpmc_send('1',x"3D44",x"0900");
    gpmc_send('1',x"3D45",x"0036");
    gpmc_send('1',x"3D46",x"0A00");
    gpmc_send('1',x"3D47",x"0035");
    gpmc_send('1',x"3D48",x"0B00");
    gpmc_send('1',x"3D49",x"0034");
    gpmc_send('1',x"3D4A",x"0C00");
    gpmc_send('1',x"3D4B",x"0033");
    gpmc_send('1',x"3D4C",x"0D00");
    gpmc_send('1',x"3D4D",x"0032");
    gpmc_send('1',x"3D4E",x"0E00");
    gpmc_send('1',x"3D4F",x"0031");
    gpmc_send('1',x"3D50",x"0F00");
    gpmc_send('1',x"3D51",x"0030");
    gpmc_send('1',x"3D52",x"1000");
    gpmc_send('1',x"3D53",x"002F");
    gpmc_send('1',x"3D54",x"1100");
    gpmc_send('1',x"3D55",x"002E");
    gpmc_send('1',x"3D56",x"1200");
    gpmc_send('1',x"3D57",x"002D");
    gpmc_send('1',x"3D58",x"1300");
    gpmc_send('1',x"3D59",x"002C");
    gpmc_send('1',x"3D5A",x"1400");
    gpmc_send('1',x"3D5B",x"002B");
    gpmc_send('1',x"3D5C",x"1500");
    gpmc_send('1',x"3D5D",x"002A");
    gpmc_send('1',x"3D5E",x"1600");
    gpmc_send('1',x"3D5F",x"0029");
    gpmc_send('1',x"3D60",x"1700");
    gpmc_send('1',x"3D61",x"0028");
    gpmc_send('1',x"3D62",x"1800");
    gpmc_send('1',x"3D63",x"0027");
    gpmc_send('1',x"3D64",x"1900");
    gpmc_send('1',x"3D65",x"0026");
    gpmc_send('1',x"3D66",x"1A00");
    gpmc_send('1',x"3D67",x"0025");
    gpmc_send('1',x"3D68",x"1B00");
    gpmc_send('1',x"3D69",x"0024");
    gpmc_send('1',x"3D6A",x"1C00");
    gpmc_send('1',x"3D6B",x"0023");
    gpmc_send('1',x"3D6C",x"1D00");
    gpmc_send('1',x"3D6D",x"0022");
    gpmc_send('1',x"3D6E",x"1E00");
    gpmc_send('1',x"3D6F",x"0021");
    gpmc_send('1',x"3D70",x"1F00");
    gpmc_send('1',x"3D71",x"0020");
    gpmc_send('1',x"3D72",x"2000");
    gpmc_send('1',x"3D73",x"001F");
    gpmc_send('1',x"3D74",x"2100");
    gpmc_send('1',x"3D75",x"001E");
    gpmc_send('1',x"3D76",x"2200");
    gpmc_send('1',x"3D77",x"001D");
    gpmc_send('1',x"3D78",x"2300");
    gpmc_send('1',x"3D79",x"001C");
    gpmc_send('1',x"3D7A",x"2400");
    gpmc_send('1',x"3D7B",x"001B");
    gpmc_send('1',x"3D7C",x"2500");
    gpmc_send('1',x"3D7D",x"001A");
    gpmc_send('1',x"3D7E",x"2600");
    gpmc_send('1',x"3D7F",x"0019");
    gpmc_send('1',x"3D80",x"2700");
    gpmc_send('1',x"3D81",x"0018");
    gpmc_send('1',x"3D82",x"2800");
    gpmc_send('1',x"3D83",x"0017");
    gpmc_send('1',x"3D84",x"2900");
    gpmc_send('1',x"3D85",x"0016");
    gpmc_send('1',x"3D86",x"2A00");
    gpmc_send('1',x"3D87",x"0015");
    gpmc_send('1',x"3D88",x"2B00");
    gpmc_send('1',x"3D89",x"0014");
    gpmc_send('1',x"3D8A",x"2C00");
    gpmc_send('1',x"3D8B",x"0013");
    gpmc_send('1',x"3D8C",x"2D00");
    gpmc_send('1',x"3D8D",x"0012");
    gpmc_send('1',x"3D8E",x"2E00");
    gpmc_send('1',x"3D8F",x"0011");
    gpmc_send('1',x"3D90",x"2F00");
    gpmc_send('1',x"3D91",x"0010");
    gpmc_send('1',x"3D92",x"3000");
    gpmc_send('1',x"3D93",x"000F");
    gpmc_send('1',x"3D94",x"3100");
    gpmc_send('1',x"3D95",x"000E");
    gpmc_send('1',x"3D96",x"3200");
    gpmc_send('1',x"3D97",x"000D");
    gpmc_send('1',x"3D98",x"3300");
    gpmc_send('1',x"3D99",x"000C");
    gpmc_send('1',x"3D9A",x"3400");
    gpmc_send('1',x"3D9B",x"000B");
    gpmc_send('1',x"3D9C",x"3500");
    gpmc_send('1',x"3D9D",x"000A");
    gpmc_send('1',x"3D9E",x"3600");
    gpmc_send('1',x"3D9F",x"0009");
    gpmc_send('1',x"3DA0",x"3700");
    gpmc_send('1',x"3DA1",x"0008");
    gpmc_send('1',x"3DA2",x"3800");
    gpmc_send('1',x"3DA3",x"0007");
    gpmc_send('1',x"3DA4",x"3900");
    gpmc_send('1',x"3DA5",x"0006");
    gpmc_send('1',x"3DA6",x"3A00");
    gpmc_send('1',x"3DA7",x"0005");
    gpmc_send('1',x"3DA8",x"3B00");
    gpmc_send('1',x"3DA9",x"0004");
    gpmc_send('1',x"3DAA",x"3C00");
    gpmc_send('1',x"3DAB",x"0003");
    gpmc_send('1',x"3DAC",x"3D00");
    gpmc_send('1',x"3DAD",x"0002");
    gpmc_send('1',x"3DAE",x"3E00");
    gpmc_send('1',x"3DAF",x"0001");
    gpmc_send('1',x"3DB0",x"3F00");
    gpmc_send('1',x"3DB1",x"0000");
    gpmc_send('1',x"3DB2",x"3F01");
    gpmc_send('1',x"3DB3",x"0000");
    gpmc_send('1',x"3DB4",x"3E02");
    gpmc_send('1',x"3DB5",x"0000");
    gpmc_send('1',x"3DB6",x"3D03");
    gpmc_send('1',x"3DB7",x"0000");
    gpmc_send('1',x"3DB8",x"3C04");
    gpmc_send('1',x"3DB9",x"0000");
    gpmc_send('1',x"3DBA",x"3B05");
    gpmc_send('1',x"3DBB",x"0000");
    gpmc_send('1',x"3DBC",x"3A06");
    gpmc_send('1',x"3DBD",x"0000");
    gpmc_send('1',x"3DBE",x"3907");
    gpmc_send('1',x"3DBF",x"0000");
    gpmc_send('1',x"3DC0",x"3808");
    gpmc_send('1',x"3DC1",x"0000");
    gpmc_send('1',x"3DC2",x"3709");
    gpmc_send('1',x"3DC3",x"0000");
    gpmc_send('1',x"3DC4",x"360A");
    gpmc_send('1',x"3DC5",x"0000");
    gpmc_send('1',x"3DC6",x"350B");
    gpmc_send('1',x"3DC7",x"0000");
    gpmc_send('1',x"3DC8",x"340C");
    gpmc_send('1',x"3DC9",x"0000");
    gpmc_send('1',x"3DCA",x"330D");
    gpmc_send('1',x"3DCB",x"0000");
    gpmc_send('1',x"3DCC",x"320E");
    gpmc_send('1',x"3DCD",x"0000");
    gpmc_send('1',x"3DCE",x"310F");
    gpmc_send('1',x"3DCF",x"0000");
    gpmc_send('1',x"3DD0",x"3010");
    gpmc_send('1',x"3DD1",x"0000");
    gpmc_send('1',x"3DD2",x"2F11");
    gpmc_send('1',x"3DD3",x"0000");
    gpmc_send('1',x"3DD4",x"2E12");
    gpmc_send('1',x"3DD5",x"0000");
    gpmc_send('1',x"3DD6",x"2D13");
    gpmc_send('1',x"3DD7",x"0000");
    gpmc_send('1',x"3DD8",x"2C14");
    gpmc_send('1',x"3DD9",x"0000");
    gpmc_send('1',x"3DDA",x"2B15");
    gpmc_send('1',x"3DDB",x"0000");
    gpmc_send('1',x"3DDC",x"2A16");
    gpmc_send('1',x"3DDD",x"0000");
    gpmc_send('1',x"3DDE",x"2917");
    gpmc_send('1',x"3DDF",x"0000");
    gpmc_send('1',x"3DE0",x"2818");
    gpmc_send('1',x"3DE1",x"0000");
    gpmc_send('1',x"3DE2",x"2719");
    gpmc_send('1',x"3DE3",x"0000");
    gpmc_send('1',x"3DE4",x"261A");
    gpmc_send('1',x"3DE5",x"0000");
    gpmc_send('1',x"3DE6",x"251B");
    gpmc_send('1',x"3DE7",x"0000");
    gpmc_send('1',x"3DE8",x"241C");
    gpmc_send('1',x"3DE9",x"0000");
    gpmc_send('1',x"3DEA",x"231D");
    gpmc_send('1',x"3DEB",x"0000");
    gpmc_send('1',x"3DEC",x"221E");
    gpmc_send('1',x"3DED",x"0000");
    gpmc_send('1',x"3DEE",x"211F");
    gpmc_send('1',x"3DEF",x"0000");
    gpmc_send('1',x"3DF0",x"2020");
    gpmc_send('1',x"3DF1",x"0000");
    gpmc_send('1',x"3DF2",x"1F21");
    gpmc_send('1',x"3DF3",x"0000");
    gpmc_send('1',x"3DF4",x"1E22");
    gpmc_send('1',x"3DF5",x"0000");
    gpmc_send('1',x"3DF6",x"1D23");
    gpmc_send('1',x"3DF7",x"0000");
    gpmc_send('1',x"3DF8",x"1C24");
    gpmc_send('1',x"3DF9",x"0000");
    gpmc_send('1',x"3DFA",x"1B25");
    gpmc_send('1',x"3DFB",x"0000");
    gpmc_send('1',x"3DFC",x"1A26");
    gpmc_send('1',x"3DFD",x"0000");
    gpmc_send('1',x"3DFE",x"1927");
    gpmc_send('1',x"3DFF",x"0000");
    gpmc_send('1',x"3E00",x"1828");
    gpmc_send('1',x"3E01",x"0000");
    gpmc_send('1',x"3E02",x"1729");
    gpmc_send('1',x"3E03",x"0000");
    gpmc_send('1',x"3E04",x"162A");
    gpmc_send('1',x"3E05",x"0000");
    gpmc_send('1',x"3E06",x"152B");
    gpmc_send('1',x"3E07",x"0000");
    gpmc_send('1',x"3E08",x"142C");
    gpmc_send('1',x"3E09",x"0000");
    gpmc_send('1',x"3E0A",x"132D");
    gpmc_send('1',x"3E0B",x"0000");
    gpmc_send('1',x"3E0C",x"122E");
    gpmc_send('1',x"3E0D",x"0000");
    gpmc_send('1',x"3E0E",x"112F");
    gpmc_send('1',x"3E0F",x"0000");
    gpmc_send('1',x"3E10",x"1030");
    gpmc_send('1',x"3E11",x"0000");
    gpmc_send('1',x"3E12",x"0F31");
    gpmc_send('1',x"3E13",x"0000");
    gpmc_send('1',x"3E14",x"0E32");
    gpmc_send('1',x"3E15",x"0000");
    gpmc_send('1',x"3E16",x"0D33");
    gpmc_send('1',x"3E17",x"0000");
    gpmc_send('1',x"3E18",x"0C34");
    gpmc_send('1',x"3E19",x"0000");
    gpmc_send('1',x"3E1A",x"0B35");
    gpmc_send('1',x"3E1B",x"0000");
    gpmc_send('1',x"3E1C",x"0A36");
    gpmc_send('1',x"3E1D",x"0000");
    gpmc_send('1',x"3E1E",x"0937");
    gpmc_send('1',x"3E1F",x"0000");
    gpmc_send('1',x"3E20",x"0838");
    gpmc_send('1',x"3E21",x"0000");
    gpmc_send('1',x"3E22",x"0739");
    gpmc_send('1',x"3E23",x"0000");
    gpmc_send('1',x"3E24",x"063A");
    gpmc_send('1',x"3E25",x"0000");
    gpmc_send('1',x"3E26",x"053B");
    gpmc_send('1',x"3E27",x"0000");
    gpmc_send('1',x"3E28",x"043C");
    gpmc_send('1',x"3E29",x"0000");
    gpmc_send('1',x"3E2A",x"033D");
    gpmc_send('1',x"3E2B",x"0000");
    gpmc_send('1',x"3E2C",x"023E");
    gpmc_send('1',x"3E2D",x"0000");
    gpmc_send('1',x"3E2E",x"013F");
    gpmc_send('1',x"3E2F",x"0000");
    gpmc_send('1',x"3E30",x"003F");
    gpmc_send('1',x"3E31",x"0000");
    gpmc_send('1',x"3E32",x"003E");
    gpmc_send('1',x"3E33",x"0001");
    gpmc_send('1',x"3E34",x"003D");
    gpmc_send('1',x"3E35",x"0002");
    gpmc_send('1',x"3E36",x"003C");
    gpmc_send('1',x"3E37",x"0003");
    gpmc_send('1',x"3E38",x"003B");
    gpmc_send('1',x"3E39",x"0004");
    gpmc_send('1',x"3E3A",x"003A");
    gpmc_send('1',x"3E3B",x"0005");
    gpmc_send('1',x"3E3C",x"0039");
    gpmc_send('1',x"3E3D",x"0006");
    gpmc_send('1',x"3E3E",x"0038");
    gpmc_send('1',x"3E3F",x"0007");
    gpmc_send('1',x"3E40",x"0037");
    gpmc_send('1',x"3E41",x"0008");
    gpmc_send('1',x"3E42",x"0036");
    gpmc_send('1',x"3E43",x"0009");
    gpmc_send('1',x"3E44",x"0035");
    gpmc_send('1',x"3E45",x"000A");
    gpmc_send('1',x"3E46",x"0034");
    gpmc_send('1',x"3E47",x"000B");
    gpmc_send('1',x"3E48",x"0033");
    gpmc_send('1',x"3E49",x"000C");
    gpmc_send('1',x"3E4A",x"0032");
    gpmc_send('1',x"3E4B",x"000D");
    gpmc_send('1',x"3E4C",x"0031");
    gpmc_send('1',x"3E4D",x"000E");
    gpmc_send('1',x"3E4E",x"0030");
    gpmc_send('1',x"3E4F",x"000F");
    gpmc_send('1',x"3E50",x"002F");
    gpmc_send('1',x"3E51",x"0010");
    gpmc_send('1',x"3E52",x"002E");
    gpmc_send('1',x"3E53",x"0011");
    gpmc_send('1',x"3E54",x"002D");
    gpmc_send('1',x"3E55",x"0012");
    gpmc_send('1',x"3E56",x"002C");
    gpmc_send('1',x"3E57",x"0013");
    gpmc_send('1',x"3E58",x"002B");
    gpmc_send('1',x"3E59",x"0014");
    gpmc_send('1',x"3E5A",x"002A");
    gpmc_send('1',x"3E5B",x"0015");
    gpmc_send('1',x"3E5C",x"0029");
    gpmc_send('1',x"3E5D",x"0016");
    gpmc_send('1',x"3E5E",x"0028");
    gpmc_send('1',x"3E5F",x"0017");
    gpmc_send('1',x"3E60",x"0027");
    gpmc_send('1',x"3E61",x"0018");
    gpmc_send('1',x"3E62",x"0026");
    gpmc_send('1',x"3E63",x"0019");
    gpmc_send('1',x"3E64",x"0025");
    gpmc_send('1',x"3E65",x"001A");
    gpmc_send('1',x"3E66",x"0024");
    gpmc_send('1',x"3E67",x"001B");
    gpmc_send('1',x"3E68",x"0023");
    gpmc_send('1',x"3E69",x"001C");
    gpmc_send('1',x"3E6A",x"0022");
    gpmc_send('1',x"3E6B",x"001D");
    gpmc_send('1',x"3E6C",x"0021");
    gpmc_send('1',x"3E6D",x"001E");
    gpmc_send('1',x"3E6E",x"0020");
    gpmc_send('1',x"3E6F",x"001F");
    gpmc_send('1',x"3E70",x"001F");
    gpmc_send('1',x"3E71",x"0020");
    gpmc_send('1',x"3E72",x"001E");
    gpmc_send('1',x"3E73",x"0021");
    gpmc_send('1',x"3E74",x"001D");
    gpmc_send('1',x"3E75",x"0022");
    gpmc_send('1',x"3E76",x"001C");
    gpmc_send('1',x"3E77",x"0023");
    gpmc_send('1',x"3E78",x"001B");
    gpmc_send('1',x"3E79",x"0024");
    gpmc_send('1',x"3E7A",x"001A");
    gpmc_send('1',x"3E7B",x"0025");
    gpmc_send('1',x"3E7C",x"0019");
    gpmc_send('1',x"3E7D",x"0026");
    gpmc_send('1',x"3E7E",x"0018");
    gpmc_send('1',x"3E7F",x"0027");
    gpmc_send('1',x"3E80",x"0017");
    gpmc_send('1',x"3E81",x"0028");
    gpmc_send('1',x"3E82",x"0016");
    gpmc_send('1',x"3E83",x"0029");
    gpmc_send('1',x"3E84",x"0015");
    gpmc_send('1',x"3E85",x"002A");
    gpmc_send('1',x"3E86",x"0014");
    gpmc_send('1',x"3E87",x"002B");
    gpmc_send('1',x"3E88",x"0013");
    gpmc_send('1',x"3E89",x"002C");
    gpmc_send('1',x"3E8A",x"0012");
    gpmc_send('1',x"3E8B",x"002D");
    gpmc_send('1',x"3E8C",x"0011");
    gpmc_send('1',x"3E8D",x"002E");
    gpmc_send('1',x"3E8E",x"0010");
    gpmc_send('1',x"3E8F",x"002F");
    gpmc_send('1',x"3E90",x"000F");
    gpmc_send('1',x"3E91",x"0030");
    gpmc_send('1',x"3E92",x"000E");
    gpmc_send('1',x"3E93",x"0031");
    gpmc_send('1',x"3E94",x"000D");
    gpmc_send('1',x"3E95",x"0032");
    gpmc_send('1',x"3E96",x"000C");
    gpmc_send('1',x"3E97",x"0033");
    gpmc_send('1',x"3E98",x"000B");
    gpmc_send('1',x"3E99",x"0034");
    gpmc_send('1',x"3E9A",x"000A");
    gpmc_send('1',x"3E9B",x"0035");
    gpmc_send('1',x"3E9C",x"0009");
    gpmc_send('1',x"3E9D",x"0036");
    gpmc_send('1',x"3E9E",x"0008");
    gpmc_send('1',x"3E9F",x"0037");
    gpmc_send('1',x"3EA0",x"0007");
    gpmc_send('1',x"3EA1",x"0038");
    gpmc_send('1',x"3EA2",x"0006");
    gpmc_send('1',x"3EA3",x"0039");
    gpmc_send('1',x"3EA4",x"0005");
    gpmc_send('1',x"3EA5",x"003A");
    gpmc_send('1',x"3EA6",x"0004");
    gpmc_send('1',x"3EA7",x"003B");
    gpmc_send('1',x"3EA8",x"0003");
    gpmc_send('1',x"3EA9",x"003C");
    gpmc_send('1',x"3EAA",x"0002");
    gpmc_send('1',x"3EAB",x"003D");
    gpmc_send('1',x"3EAC",x"0001");
    gpmc_send('1',x"3EAD",x"003E");
    gpmc_send('1',x"3EAE",x"0000");
    gpmc_send('1',x"3EAF",x"003F");
    gpmc_send('1',x"3EB0",x"0100");
    gpmc_send('1',x"3EB1",x"003E");
    gpmc_send('1',x"3EB2",x"0200");
    gpmc_send('1',x"3EB3",x"003D");
    gpmc_send('1',x"3EB4",x"0300");
    gpmc_send('1',x"3EB5",x"003C");
    gpmc_send('1',x"3EB6",x"0400");
    gpmc_send('1',x"3EB7",x"003B");
    gpmc_send('1',x"3EB8",x"0500");
    gpmc_send('1',x"3EB9",x"003A");
    gpmc_send('1',x"3EBA",x"0600");
    gpmc_send('1',x"3EBB",x"0039");
    gpmc_send('1',x"3EBC",x"0700");
    gpmc_send('1',x"3EBD",x"0038");
    gpmc_send('1',x"3EBE",x"0800");
    gpmc_send('1',x"3EBF",x"0037");
    gpmc_send('1',x"3EC0",x"0900");
    gpmc_send('1',x"3EC1",x"0036");
    gpmc_send('1',x"3EC2",x"0A00");
    gpmc_send('1',x"3EC3",x"0035");
    gpmc_send('1',x"3EC4",x"0B00");
    gpmc_send('1',x"3EC5",x"0034");
    gpmc_send('1',x"3EC6",x"0C00");
    gpmc_send('1',x"3EC7",x"0033");
    gpmc_send('1',x"3EC8",x"0D00");
    gpmc_send('1',x"3EC9",x"0032");
    gpmc_send('1',x"3ECA",x"0E00");
    gpmc_send('1',x"3ECB",x"0031");
    gpmc_send('1',x"3ECC",x"0F00");
    gpmc_send('1',x"3ECD",x"0030");
    gpmc_send('1',x"3ECE",x"1000");
    gpmc_send('1',x"3ECF",x"002F");
    gpmc_send('1',x"3ED0",x"1100");
    gpmc_send('1',x"3ED1",x"002E");
    gpmc_send('1',x"3ED2",x"1200");
    gpmc_send('1',x"3ED3",x"002D");
    gpmc_send('1',x"3ED4",x"1300");
    gpmc_send('1',x"3ED5",x"002C");
    gpmc_send('1',x"3ED6",x"1400");
    gpmc_send('1',x"3ED7",x"002B");
    gpmc_send('1',x"3ED8",x"1500");
    gpmc_send('1',x"3ED9",x"002A");
    gpmc_send('1',x"3EDA",x"1600");
    gpmc_send('1',x"3EDB",x"0029");
    gpmc_send('1',x"3EDC",x"1700");
    gpmc_send('1',x"3EDD",x"0028");
    gpmc_send('1',x"3EDE",x"1800");
    gpmc_send('1',x"3EDF",x"0027");
    gpmc_send('1',x"3EE0",x"1900");
    gpmc_send('1',x"3EE1",x"0026");
    gpmc_send('1',x"3EE2",x"1A00");
    gpmc_send('1',x"3EE3",x"0025");
    gpmc_send('1',x"3EE4",x"1B00");
    gpmc_send('1',x"3EE5",x"0024");
    gpmc_send('1',x"3EE6",x"1C00");
    gpmc_send('1',x"3EE7",x"0023");
    gpmc_send('1',x"3EE8",x"1D00");
    gpmc_send('1',x"3EE9",x"0022");
    gpmc_send('1',x"3EEA",x"1E00");
    gpmc_send('1',x"3EEB",x"0021");
    gpmc_send('1',x"3EEC",x"1F00");
    gpmc_send('1',x"3EED",x"0020");
    gpmc_send('1',x"3EEE",x"2000");
    gpmc_send('1',x"3EEF",x"001F");
    gpmc_send('1',x"3EF0",x"2100");
    gpmc_send('1',x"3EF1",x"001E");
    gpmc_send('1',x"3EF2",x"2200");
    gpmc_send('1',x"3EF3",x"001D");
    gpmc_send('1',x"3EF4",x"2300");
    gpmc_send('1',x"3EF5",x"001C");
    gpmc_send('1',x"3EF6",x"2400");
    gpmc_send('1',x"3EF7",x"001B");
    gpmc_send('1',x"3EF8",x"2500");
    gpmc_send('1',x"3EF9",x"001A");
    gpmc_send('1',x"3EFA",x"2600");
    gpmc_send('1',x"3EFB",x"0019");
    gpmc_send('1',x"3EFC",x"2700");
    gpmc_send('1',x"3EFD",x"0018");
    gpmc_send('1',x"3EFE",x"2800");
    gpmc_send('1',x"3EFF",x"0017");
    gpmc_send('1',x"3F00",x"2900");
    gpmc_send('1',x"3F01",x"0016");
    gpmc_send('1',x"3F02",x"2A00");
    gpmc_send('1',x"3F03",x"0015");
    gpmc_send('1',x"3F04",x"2B00");
    gpmc_send('1',x"3F05",x"0014");
    gpmc_send('1',x"3F06",x"2C00");
    gpmc_send('1',x"3F07",x"0013");
    gpmc_send('1',x"3F08",x"2D00");
    gpmc_send('1',x"3F09",x"0012");
    gpmc_send('1',x"3F0A",x"2E00");
    gpmc_send('1',x"3F0B",x"0011");
    gpmc_send('1',x"3F0C",x"2F00");
    gpmc_send('1',x"3F0D",x"0010");
    gpmc_send('1',x"3F0E",x"3000");
    gpmc_send('1',x"3F0F",x"000F");
    gpmc_send('1',x"3F10",x"3100");
    gpmc_send('1',x"3F11",x"000E");
    gpmc_send('1',x"3F12",x"3200");
    gpmc_send('1',x"3F13",x"000D");
    gpmc_send('1',x"3F14",x"3300");
    gpmc_send('1',x"3F15",x"000C");
    gpmc_send('1',x"3F16",x"3400");
    gpmc_send('1',x"3F17",x"000B");
    gpmc_send('1',x"3F18",x"3500");
    gpmc_send('1',x"3F19",x"000A");
    gpmc_send('1',x"3F1A",x"3600");
    gpmc_send('1',x"3F1B",x"0009");
    gpmc_send('1',x"3F1C",x"3700");
    gpmc_send('1',x"3F1D",x"0008");
    gpmc_send('1',x"3F1E",x"3800");
    gpmc_send('1',x"3F1F",x"0007");
    gpmc_send('1',x"3F20",x"3900");
    gpmc_send('1',x"3F21",x"0006");
    gpmc_send('1',x"3F22",x"3A00");
    gpmc_send('1',x"3F23",x"0005");
    gpmc_send('1',x"3F24",x"3B00");
    gpmc_send('1',x"3F25",x"0004");
    gpmc_send('1',x"3F26",x"3C00");
    gpmc_send('1',x"3F27",x"0003");
    gpmc_send('1',x"3F28",x"3D00");
    gpmc_send('1',x"3F29",x"0002");
    gpmc_send('1',x"3F2A",x"3E00");
    gpmc_send('1',x"3F2B",x"0001");
    gpmc_send('1',x"3F2C",x"3F00");
    gpmc_send('1',x"3F2D",x"0000");
    gpmc_send('1',x"3F2E",x"3F01");
    gpmc_send('1',x"3F2F",x"0000");
    gpmc_send('1',x"3F30",x"3E02");
    gpmc_send('1',x"3F31",x"0000");
    gpmc_send('1',x"3F32",x"3D03");
    gpmc_send('1',x"3F33",x"0000");
    gpmc_send('1',x"3F34",x"3C04");
    gpmc_send('1',x"3F35",x"0000");
    gpmc_send('1',x"3F36",x"3B05");
    gpmc_send('1',x"3F37",x"0000");
    gpmc_send('1',x"3F38",x"3A06");
    gpmc_send('1',x"3F39",x"0000");
    gpmc_send('1',x"3F3A",x"3907");
    gpmc_send('1',x"3F3B",x"0000");
    gpmc_send('1',x"3F3C",x"3808");
    gpmc_send('1',x"3F3D",x"0000");
    gpmc_send('1',x"3F3E",x"3709");
    gpmc_send('1',x"3F3F",x"0000");
    gpmc_send('1',x"3F40",x"360A");
    gpmc_send('1',x"3F41",x"0000");
    gpmc_send('1',x"3F42",x"350B");
    gpmc_send('1',x"3F43",x"0000");
    gpmc_send('1',x"3F44",x"340C");
    gpmc_send('1',x"3F45",x"0000");
    gpmc_send('1',x"3F46",x"330D");
    gpmc_send('1',x"3F47",x"0000");
    gpmc_send('1',x"3F48",x"320E");
    gpmc_send('1',x"3F49",x"0000");
    gpmc_send('1',x"3F4A",x"310F");
    gpmc_send('1',x"3F4B",x"0000");
    gpmc_send('1',x"3F4C",x"3010");
    gpmc_send('1',x"3F4D",x"0000");
    gpmc_send('1',x"3F4E",x"2F11");
    gpmc_send('1',x"3F4F",x"0000");
    gpmc_send('1',x"3F50",x"2E12");
    gpmc_send('1',x"3F51",x"0000");
    gpmc_send('1',x"3F52",x"2D13");
    gpmc_send('1',x"3F53",x"0000");
    gpmc_send('1',x"3F54",x"2C14");
    gpmc_send('1',x"3F55",x"0000");
    gpmc_send('1',x"3F56",x"2B15");
    gpmc_send('1',x"3F57",x"0000");
    gpmc_send('1',x"3F58",x"2A16");
    gpmc_send('1',x"3F59",x"0000");
    gpmc_send('1',x"3F5A",x"2917");
    gpmc_send('1',x"3F5B",x"0000");
    gpmc_send('1',x"3F5C",x"2818");
    gpmc_send('1',x"3F5D",x"0000");
    gpmc_send('1',x"3F5E",x"2719");
    gpmc_send('1',x"3F5F",x"0000");
    gpmc_send('1',x"3F60",x"261A");
    gpmc_send('1',x"3F61",x"0000");
    gpmc_send('1',x"3F62",x"251B");
    gpmc_send('1',x"3F63",x"0000");
    gpmc_send('1',x"3F64",x"241C");
    gpmc_send('1',x"3F65",x"0000");
    gpmc_send('1',x"3F66",x"231D");
    gpmc_send('1',x"3F67",x"0000");
    gpmc_send('1',x"3F68",x"221E");
    gpmc_send('1',x"3F69",x"0000");
    gpmc_send('1',x"3F6A",x"211F");
    gpmc_send('1',x"3F6B",x"0000");
    gpmc_send('1',x"3F6C",x"2020");
    gpmc_send('1',x"3F6D",x"0000");
    gpmc_send('1',x"3F6E",x"1F21");
    gpmc_send('1',x"3F6F",x"0000");
    gpmc_send('1',x"3F70",x"1E22");
    gpmc_send('1',x"3F71",x"0000");
    gpmc_send('1',x"3F72",x"1D23");
    gpmc_send('1',x"3F73",x"0000");
    gpmc_send('1',x"3F74",x"1C24");
    gpmc_send('1',x"3F75",x"0000");
    gpmc_send('1',x"3F76",x"1B25");
    gpmc_send('1',x"3F77",x"0000");
    gpmc_send('1',x"3F78",x"1A26");
    gpmc_send('1',x"3F79",x"0000");
    gpmc_send('1',x"3F7A",x"1927");
    gpmc_send('1',x"3F7B",x"0000");
    gpmc_send('1',x"3F7C",x"1828");
    gpmc_send('1',x"3F7D",x"0000");
    gpmc_send('1',x"3F7E",x"1729");
    gpmc_send('1',x"3F7F",x"0000");
    gpmc_send('1',x"3F80",x"162A");
    gpmc_send('1',x"3F81",x"0000");
    gpmc_send('1',x"3F82",x"152B");
    gpmc_send('1',x"3F83",x"0000");
    gpmc_send('1',x"3F84",x"142C");
    gpmc_send('1',x"3F85",x"0000");
    gpmc_send('1',x"3F86",x"132D");
    gpmc_send('1',x"3F87",x"0000");
    gpmc_send('1',x"3F88",x"122E");
    gpmc_send('1',x"3F89",x"0000");
    gpmc_send('1',x"3F8A",x"112F");
    gpmc_send('1',x"3F8B",x"0000");
    gpmc_send('1',x"3F8C",x"1030");
    gpmc_send('1',x"3F8D",x"0000");
    gpmc_send('1',x"3F8E",x"0F31");
    gpmc_send('1',x"3F8F",x"0000");
    gpmc_send('1',x"3F90",x"0E32");
    gpmc_send('1',x"3F91",x"0000");
    gpmc_send('1',x"3F92",x"0D33");
    gpmc_send('1',x"3F93",x"0000");
    gpmc_send('1',x"3F94",x"0C34");
    gpmc_send('1',x"3F95",x"0000");
    gpmc_send('1',x"3F96",x"0B35");
    gpmc_send('1',x"3F97",x"0000");
    gpmc_send('1',x"3F98",x"0A36");
    gpmc_send('1',x"3F99",x"0000");
    gpmc_send('1',x"3F9A",x"0937");
    gpmc_send('1',x"3F9B",x"0000");
    gpmc_send('1',x"3F9C",x"0838");
    gpmc_send('1',x"3F9D",x"0000");
    gpmc_send('1',x"3F9E",x"0739");
    gpmc_send('1',x"3F9F",x"0000");
    gpmc_send('1',x"3FA0",x"063A");
    gpmc_send('1',x"3FA1",x"0000");
    gpmc_send('1',x"3FA2",x"053B");
    gpmc_send('1',x"3FA3",x"0000");
    gpmc_send('1',x"3FA4",x"043C");
    gpmc_send('1',x"3FA5",x"0000");
    gpmc_send('1',x"3FA6",x"033D");
    gpmc_send('1',x"3FA7",x"0000");
    gpmc_send('1',x"3FA8",x"023E");
    gpmc_send('1',x"3FA9",x"0000");
    gpmc_send('1',x"3FAA",x"013F");
    gpmc_send('1',x"3FAB",x"0000");
    gpmc_send('1',x"3FAC",x"003F");
    gpmc_send('1',x"3FAD",x"0000");
    gpmc_send('1',x"3FAE",x"003E");
    gpmc_send('1',x"3FAF",x"0001");
    gpmc_send('1',x"3FB0",x"003D");
    gpmc_send('1',x"3FB1",x"0002");
    gpmc_send('1',x"3FB2",x"003C");
    gpmc_send('1',x"3FB3",x"0003");
    gpmc_send('1',x"3FB4",x"003B");
    gpmc_send('1',x"3FB5",x"0004");
    gpmc_send('1',x"3FB6",x"003A");
    gpmc_send('1',x"3FB7",x"0005");
    gpmc_send('1',x"3FB8",x"0039");
    gpmc_send('1',x"3FB9",x"0006");
    gpmc_send('1',x"3FBA",x"0038");
    gpmc_send('1',x"3FBB",x"0007");
    gpmc_send('1',x"3FBC",x"0037");
    gpmc_send('1',x"3FBD",x"0008");
    gpmc_send('1',x"3FBE",x"0036");
    gpmc_send('1',x"3FBF",x"0009");
    gpmc_send('1',x"3FC0",x"0035");
    gpmc_send('1',x"3FC1",x"000A");
    gpmc_send('1',x"3FC2",x"0034");
    gpmc_send('1',x"3FC3",x"000B");
    gpmc_send('1',x"3FC4",x"0033");
    gpmc_send('1',x"3FC5",x"000C");
    gpmc_send('1',x"3FC6",x"0032");
    gpmc_send('1',x"3FC7",x"000D");
    gpmc_send('1',x"3FC8",x"0031");
    gpmc_send('1',x"3FC9",x"000E");
    gpmc_send('1',x"3FCA",x"0030");
    gpmc_send('1',x"3FCB",x"000F");
    gpmc_send('1',x"3FCC",x"002F");
    gpmc_send('1',x"3FCD",x"0010");
    gpmc_send('1',x"3FCE",x"002E");
    gpmc_send('1',x"3FCF",x"0011");
    gpmc_send('1',x"3FD0",x"002D");
    gpmc_send('1',x"3FD1",x"0012");
    gpmc_send('1',x"3FD2",x"002C");
    gpmc_send('1',x"3FD3",x"0013");
    gpmc_send('1',x"3FD4",x"002B");
    gpmc_send('1',x"3FD5",x"0014");
    gpmc_send('1',x"3FD6",x"002A");
    gpmc_send('1',x"3FD7",x"0015");
    gpmc_send('1',x"3FD8",x"0029");
    gpmc_send('1',x"3FD9",x"0016");
    gpmc_send('1',x"3FDA",x"0028");
    gpmc_send('1',x"3FDB",x"0017");
    gpmc_send('1',x"3FDC",x"0027");
    gpmc_send('1',x"3FDD",x"0018");
    gpmc_send('1',x"3FDE",x"0026");
    gpmc_send('1',x"3FDF",x"0019");
    gpmc_send('1',x"3FE0",x"0025");
    gpmc_send('1',x"3FE1",x"001A");
    gpmc_send('1',x"3FE2",x"0024");
    gpmc_send('1',x"3FE3",x"001B");
    gpmc_send('1',x"3FE4",x"0023");
    gpmc_send('1',x"3FE5",x"001C");
    gpmc_send('1',x"3FE6",x"0022");
    gpmc_send('1',x"3FE7",x"001D");
    gpmc_send('1',x"3FE8",x"0021");
    gpmc_send('1',x"3FE9",x"001E");
    gpmc_send('1',x"3FEA",x"0020");
    gpmc_send('1',x"3FEB",x"001F");
    gpmc_send('1',x"3FEC",x"001F");
    gpmc_send('1',x"3FED",x"0020");
    gpmc_send('1',x"3FEE",x"001E");
    gpmc_send('1',x"3FEF",x"0021");
    gpmc_send('1',x"3FF0",x"001D");
    gpmc_send('1',x"3FF1",x"0022");
    gpmc_send('1',x"3FF2",x"001C");
    gpmc_send('1',x"3FF3",x"0023");
    gpmc_send('1',x"3FF4",x"001B");
    gpmc_send('1',x"3FF5",x"0024");
    gpmc_send('1',x"3FF6",x"001A");
    gpmc_send('1',x"3FF7",x"0025");
    gpmc_send('1',x"3FF8",x"0019");
    gpmc_send('1',x"3FF9",x"0026");
    gpmc_send('1',x"3FFA",x"0018");
    gpmc_send('1',x"3FFB",x"0027");
    gpmc_send('1',x"3FFC",x"0017");
    gpmc_send('1',x"3FFD",x"0028");

    wait;
    end process;

end architecture;